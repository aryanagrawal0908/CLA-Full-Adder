magic
tech scmos
timestamp 1731333225
<< nwell >>
rect 241 202 273 328
rect 293 202 325 328
rect 345 264 377 328
rect 397 264 429 328
rect 442 272 506 336
<< ntransistor >>
rect 457 241 459 261
rect 489 241 491 261
rect 360 217 362 237
rect 412 217 414 237
rect 256 170 258 190
rect 308 170 310 190
rect 360 170 362 190
rect 412 170 414 190
<< ptransistor >>
rect 256 273 258 313
rect 308 273 310 313
rect 360 273 362 313
rect 412 273 414 313
rect 457 281 459 321
rect 489 281 491 321
rect 256 211 258 251
rect 308 211 310 251
<< ndiffusion >>
rect 456 241 457 261
rect 459 241 460 261
rect 488 241 489 261
rect 491 241 492 261
rect 359 217 360 237
rect 362 217 363 237
rect 411 217 412 237
rect 414 217 415 237
rect 255 170 256 190
rect 258 170 259 190
rect 307 170 308 190
rect 310 170 311 190
rect 359 170 360 190
rect 362 170 363 190
rect 411 170 412 190
rect 414 170 415 190
<< pdiffusion >>
rect 255 273 256 313
rect 258 273 259 313
rect 307 273 308 313
rect 310 273 311 313
rect 359 273 360 313
rect 362 273 363 313
rect 411 273 412 313
rect 414 273 415 313
rect 456 281 457 321
rect 459 281 460 321
rect 488 281 489 321
rect 491 281 492 321
rect 255 211 256 251
rect 258 211 259 251
rect 307 211 308 251
rect 310 211 311 251
<< ndcontact >>
rect 452 241 456 261
rect 460 241 464 261
rect 484 241 488 261
rect 492 241 496 261
rect 355 217 359 237
rect 363 217 367 237
rect 407 217 411 237
rect 415 217 419 237
rect 251 170 255 190
rect 259 170 263 190
rect 303 170 307 190
rect 311 170 315 190
rect 355 170 359 190
rect 363 170 367 190
rect 407 170 411 190
rect 415 170 419 190
<< pdcontact >>
rect 251 273 255 313
rect 259 273 263 313
rect 303 273 307 313
rect 311 273 315 313
rect 355 273 359 313
rect 363 273 367 313
rect 407 273 411 313
rect 415 273 419 313
rect 452 281 456 321
rect 460 281 464 321
rect 484 281 488 321
rect 492 281 496 321
rect 251 211 255 251
rect 259 211 263 251
rect 303 211 307 251
rect 311 211 315 251
<< psubstratepcontact >>
rect 444 228 448 232
rect 468 228 472 232
rect 476 228 480 232
rect 500 228 504 232
rect 268 157 272 161
rect 320 157 324 161
rect 372 157 376 161
rect 424 157 428 161
<< nsubstratencontact >>
rect 445 329 449 333
rect 467 329 471 333
rect 477 329 481 333
rect 499 329 503 333
rect 244 321 248 325
rect 266 321 270 325
rect 296 321 300 325
rect 318 321 322 325
rect 348 321 352 325
rect 370 321 374 325
rect 400 321 404 325
rect 422 321 426 325
<< polysilicon >>
rect 457 321 459 325
rect 489 321 491 325
rect 256 313 258 317
rect 308 313 310 317
rect 360 313 362 317
rect 412 313 414 317
rect 256 264 258 273
rect 308 264 310 273
rect 360 264 362 273
rect 412 264 414 273
rect 457 261 459 281
rect 489 261 491 281
rect 256 251 258 255
rect 308 251 310 255
rect 360 237 362 246
rect 412 237 414 246
rect 457 237 459 241
rect 489 237 491 241
rect 360 214 362 217
rect 412 214 414 217
rect 256 202 258 211
rect 308 202 310 211
rect 256 190 258 198
rect 308 190 310 198
rect 360 190 362 198
rect 412 190 414 198
rect 256 166 258 170
rect 308 166 310 170
rect 360 166 362 170
rect 412 166 414 170
<< polycontact >>
rect 251 264 256 269
rect 303 264 308 269
rect 355 264 360 269
rect 407 264 412 269
rect 452 264 457 269
rect 484 264 489 269
rect 355 241 360 246
rect 407 241 412 246
rect 251 202 256 207
rect 303 202 308 207
rect 251 193 256 198
rect 303 193 308 198
rect 355 193 360 198
rect 407 193 412 198
<< metal1 >>
rect 442 333 506 336
rect 442 329 445 333
rect 449 329 467 333
rect 471 329 477 333
rect 481 329 499 333
rect 503 329 506 333
rect 241 325 429 328
rect 442 327 506 329
rect 241 321 244 325
rect 248 321 266 325
rect 270 321 296 325
rect 300 321 318 325
rect 322 321 348 325
rect 352 321 370 325
rect 374 321 400 325
rect 404 321 422 325
rect 426 321 429 325
rect 241 319 429 321
rect 452 321 456 327
rect 484 321 488 327
rect 251 313 255 319
rect 303 313 307 319
rect 355 313 359 319
rect 407 313 411 319
rect 228 264 251 269
rect 228 198 233 264
rect 259 260 263 273
rect 251 256 263 260
rect 281 264 303 269
rect 251 251 255 256
rect 246 202 251 207
rect 259 198 263 211
rect 281 198 286 264
rect 311 260 315 273
rect 363 269 367 273
rect 415 269 419 273
rect 460 269 464 281
rect 492 269 496 281
rect 303 256 315 260
rect 333 264 355 269
rect 363 264 407 269
rect 415 264 452 269
rect 460 264 484 269
rect 492 264 506 269
rect 303 251 307 256
rect 298 202 303 207
rect 311 198 315 211
rect 333 198 338 264
rect 352 241 355 246
rect 363 237 367 264
rect 355 206 359 217
rect 355 202 367 206
rect 228 193 251 198
rect 259 193 303 198
rect 311 193 355 198
rect 259 190 263 193
rect 311 190 315 193
rect 363 190 367 202
rect 385 198 390 264
rect 404 241 407 246
rect 415 237 419 264
rect 460 261 464 264
rect 492 261 496 264
rect 452 234 456 241
rect 484 234 488 241
rect 442 232 506 234
rect 442 228 444 232
rect 448 228 468 232
rect 472 228 476 232
rect 480 228 500 232
rect 504 228 506 232
rect 442 226 506 228
rect 407 206 411 217
rect 407 202 419 206
rect 385 193 407 198
rect 415 190 419 202
rect 251 162 255 170
rect 303 162 307 170
rect 355 162 359 170
rect 407 162 411 170
rect 241 161 429 162
rect 241 157 268 161
rect 272 157 320 161
rect 324 157 372 161
rect 376 157 424 161
rect 428 157 429 161
rect 241 156 429 157
rect 234 143 241 148
rect 246 143 293 148
rect 298 143 347 148
rect 352 143 399 148
<< m2contact >>
rect 241 202 246 207
rect 293 202 298 207
rect 347 241 352 246
rect 399 241 404 246
rect 241 143 246 148
rect 293 143 298 148
rect 347 143 352 148
rect 399 143 404 148
<< metal2 >>
rect 241 148 246 202
rect 293 148 298 202
rect 347 148 352 241
rect 399 148 404 241
<< labels >>
rlabel metal1 257 324 257 324 5 vdd
rlabel metal1 257 159 257 159 1 gnd
rlabel metal1 309 324 309 324 5 vdd
rlabel metal1 309 159 309 159 1 gnd
rlabel metal1 361 159 361 159 1 gnd
rlabel metal1 361 324 361 324 5 vdd
rlabel metal1 413 159 413 159 1 gnd
rlabel metal1 413 324 413 324 5 vdd
rlabel metal1 230 234 230 234 1 d
rlabel metal1 489 230 489 230 1 gnd
rlabel metal1 490 332 490 332 5 vdd
rlabel metal1 457 230 457 230 1 gnd
rlabel metal1 458 332 458 332 5 vdd
rlabel metal1 236 145 236 145 1 clk
rlabel metal1 261 265 261 265 1 d1
rlabel metal1 283 235 283 235 1 a
rlabel metal1 313 266 313 266 1 d2
rlabel metal1 335 234 335 234 1 q1
rlabel metal1 365 198 365 198 1 d3
rlabel metal1 388 233 388 233 1 b
rlabel metal1 417 197 417 197 1 d4
rlabel metal1 436 266 436 266 1 qmid
rlabel metal1 471 266 471 266 1 qnot
rlabel metal1 501 267 501 267 7 q
<< end >>
