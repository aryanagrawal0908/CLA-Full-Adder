magic
tech scmos
timestamp 1731255356
<< nwell >>
rect 253 245 317 277
rect 253 194 317 226
rect 395 224 427 288
rect 133 99 165 163
rect 171 99 203 163
rect 404 107 474 171
rect 368 64 400 98
rect 489 64 553 96
rect -9 0 55 32
rect -9 -51 55 -19
rect 133 -21 165 43
rect 298 -21 368 43
rect 489 13 553 45
rect 631 43 663 107
rect 262 -64 294 -30
rect 133 -191 165 -127
rect 171 -191 203 -127
rect 481 -183 551 -119
rect 445 -226 477 -192
rect -9 -290 55 -258
rect -9 -341 55 -309
rect 133 -311 165 -247
rect 378 -311 448 -247
rect 601 -305 671 -241
rect 342 -354 374 -320
rect 565 -348 597 -314
rect 691 -348 755 -316
rect 306 -437 376 -373
rect 691 -399 755 -367
rect 833 -369 865 -305
rect 270 -480 302 -446
rect 435 -467 505 -403
rect 399 -510 431 -476
rect 133 -608 165 -544
rect 171 -608 203 -544
rect 638 -600 708 -536
rect 602 -643 634 -609
rect -9 -707 55 -675
rect -9 -758 55 -726
rect 133 -728 165 -664
rect 330 -728 400 -664
rect 805 -737 875 -673
rect 294 -771 326 -737
rect 769 -780 801 -746
rect 890 -780 954 -748
rect 330 -872 400 -808
rect 890 -831 954 -799
rect 1032 -801 1064 -737
rect 294 -915 326 -881
rect 459 -902 529 -838
rect 423 -945 455 -911
rect 634 -956 704 -892
rect 333 -1042 403 -978
rect 598 -999 630 -965
rect 297 -1085 329 -1051
rect 464 -1072 534 -1008
rect 428 -1115 460 -1081
rect 333 -1186 403 -1122
rect 297 -1229 329 -1195
rect 133 -1309 165 -1245
rect 171 -1309 203 -1245
rect -9 -1408 55 -1376
rect -9 -1459 55 -1427
rect 133 -1429 165 -1365
rect 342 -1429 412 -1365
rect 496 -1389 566 -1325
rect 460 -1432 492 -1398
rect 306 -1472 338 -1438
rect 845 -1485 915 -1421
rect 342 -1573 412 -1509
rect 809 -1528 841 -1494
rect 306 -1616 338 -1582
rect 471 -1603 541 -1539
rect 435 -1646 467 -1612
rect 605 -1664 675 -1600
rect 345 -1743 415 -1679
rect 569 -1707 601 -1673
rect 309 -1786 341 -1752
rect 476 -1773 546 -1709
rect 440 -1816 472 -1782
rect 345 -1887 415 -1823
rect 734 -1853 804 -1789
rect 698 -1896 730 -1862
rect 309 -1930 341 -1896
rect 345 -2014 415 -1950
rect 309 -2057 341 -2023
rect 476 -2044 546 -1980
rect 440 -2087 472 -2053
rect 611 -2074 681 -2010
rect 345 -2158 415 -2094
rect 575 -2117 607 -2083
rect 309 -2201 341 -2167
<< ntransistor >>
rect 328 260 348 262
rect 378 252 380 272
rect 378 220 380 240
rect 328 209 348 211
rect 410 193 412 213
rect 116 101 118 121
rect 116 69 118 89
rect 383 106 385 126
rect 148 68 150 88
rect 186 68 188 88
rect 419 76 421 96
rect 457 76 459 96
rect 564 79 584 81
rect 614 71 616 91
rect 614 39 616 59
rect 564 28 584 30
rect 66 15 86 17
rect 116 7 118 27
rect 116 -25 118 -5
rect 277 -22 279 -2
rect 646 12 648 32
rect 66 -36 86 -34
rect 148 -52 150 -32
rect 313 -52 315 -32
rect 351 -52 353 -32
rect 116 -189 118 -169
rect 116 -221 118 -201
rect 460 -184 462 -164
rect 148 -222 150 -202
rect 186 -222 188 -202
rect 496 -214 498 -194
rect 534 -214 536 -194
rect 66 -275 86 -273
rect 116 -283 118 -263
rect 116 -315 118 -295
rect 357 -312 359 -292
rect 66 -326 86 -324
rect 148 -342 150 -322
rect 580 -306 582 -286
rect 393 -342 395 -322
rect 431 -342 433 -322
rect 616 -336 618 -316
rect 654 -336 656 -316
rect 766 -333 786 -331
rect 816 -341 818 -321
rect 816 -373 818 -353
rect 766 -384 786 -382
rect 285 -438 287 -418
rect 848 -400 850 -380
rect 321 -468 323 -448
rect 359 -468 361 -448
rect 414 -468 416 -448
rect 450 -498 452 -478
rect 488 -498 490 -478
rect 116 -606 118 -586
rect 116 -638 118 -618
rect 617 -601 619 -581
rect 148 -639 150 -619
rect 186 -639 188 -619
rect 653 -631 655 -611
rect 691 -631 693 -611
rect 66 -692 86 -690
rect 116 -700 118 -680
rect 116 -732 118 -712
rect 309 -729 311 -709
rect 66 -743 86 -741
rect 148 -759 150 -739
rect 784 -738 786 -718
rect 345 -759 347 -739
rect 383 -759 385 -739
rect 820 -768 822 -748
rect 858 -768 860 -748
rect 965 -765 985 -763
rect 1015 -773 1017 -753
rect 1015 -805 1017 -785
rect 965 -816 985 -814
rect 309 -873 311 -853
rect 1047 -832 1049 -812
rect 345 -903 347 -883
rect 383 -903 385 -883
rect 438 -903 440 -883
rect 474 -933 476 -913
rect 512 -933 514 -913
rect 613 -957 615 -937
rect 649 -987 651 -967
rect 687 -987 689 -967
rect 312 -1043 314 -1023
rect 348 -1073 350 -1053
rect 386 -1073 388 -1053
rect 443 -1073 445 -1053
rect 479 -1103 481 -1083
rect 517 -1103 519 -1083
rect 312 -1187 314 -1167
rect 348 -1217 350 -1197
rect 386 -1217 388 -1197
rect 116 -1307 118 -1287
rect 116 -1339 118 -1319
rect 148 -1340 150 -1320
rect 186 -1340 188 -1320
rect 66 -1393 86 -1391
rect 116 -1401 118 -1381
rect 116 -1433 118 -1413
rect 321 -1430 323 -1410
rect 475 -1390 477 -1370
rect 66 -1444 86 -1442
rect 148 -1460 150 -1440
rect 511 -1420 513 -1400
rect 549 -1420 551 -1400
rect 357 -1460 359 -1440
rect 395 -1460 397 -1440
rect 824 -1486 826 -1466
rect 860 -1516 862 -1496
rect 898 -1516 900 -1496
rect 321 -1574 323 -1554
rect 357 -1604 359 -1584
rect 395 -1604 397 -1584
rect 450 -1604 452 -1584
rect 486 -1634 488 -1614
rect 524 -1634 526 -1614
rect 584 -1665 586 -1645
rect 324 -1744 326 -1724
rect 620 -1695 622 -1675
rect 658 -1695 660 -1675
rect 360 -1774 362 -1754
rect 398 -1774 400 -1754
rect 455 -1774 457 -1754
rect 491 -1804 493 -1784
rect 529 -1804 531 -1784
rect 324 -1888 326 -1868
rect 713 -1854 715 -1834
rect 749 -1884 751 -1864
rect 787 -1884 789 -1864
rect 360 -1918 362 -1898
rect 398 -1918 400 -1898
rect 324 -2015 326 -1995
rect 360 -2045 362 -2025
rect 398 -2045 400 -2025
rect 455 -2045 457 -2025
rect 491 -2075 493 -2055
rect 529 -2075 531 -2055
rect 590 -2075 592 -2055
rect 324 -2159 326 -2139
rect 626 -2105 628 -2085
rect 664 -2105 666 -2085
rect 360 -2189 362 -2169
rect 398 -2189 400 -2169
<< ptransistor >>
rect 268 260 308 262
rect 410 233 412 273
rect 268 209 308 211
rect 148 108 150 148
rect 186 108 188 148
rect 419 116 421 156
rect 457 116 459 156
rect 383 71 385 91
rect 504 79 544 81
rect 646 52 648 92
rect 504 28 544 30
rect 6 15 46 17
rect 148 -12 150 28
rect 313 -12 315 28
rect 351 -12 353 28
rect 6 -36 46 -34
rect 277 -57 279 -37
rect 148 -182 150 -142
rect 186 -182 188 -142
rect 496 -174 498 -134
rect 534 -174 536 -134
rect 460 -219 462 -199
rect 6 -275 46 -273
rect 148 -302 150 -262
rect 393 -302 395 -262
rect 431 -302 433 -262
rect 6 -326 46 -324
rect 616 -296 618 -256
rect 654 -296 656 -256
rect 357 -347 359 -327
rect 580 -341 582 -321
rect 706 -333 746 -331
rect 848 -360 850 -320
rect 706 -384 746 -382
rect 321 -428 323 -388
rect 359 -428 361 -388
rect 285 -473 287 -453
rect 450 -458 452 -418
rect 488 -458 490 -418
rect 414 -503 416 -483
rect 148 -599 150 -559
rect 186 -599 188 -559
rect 653 -591 655 -551
rect 691 -591 693 -551
rect 617 -636 619 -616
rect 6 -692 46 -690
rect 148 -719 150 -679
rect 345 -719 347 -679
rect 383 -719 385 -679
rect 6 -743 46 -741
rect 820 -728 822 -688
rect 858 -728 860 -688
rect 309 -764 311 -744
rect 784 -773 786 -753
rect 905 -765 945 -763
rect 1047 -792 1049 -752
rect 905 -816 945 -814
rect 345 -863 347 -823
rect 383 -863 385 -823
rect 309 -908 311 -888
rect 474 -893 476 -853
rect 512 -893 514 -853
rect 438 -938 440 -918
rect 649 -947 651 -907
rect 687 -947 689 -907
rect 613 -992 615 -972
rect 348 -1033 350 -993
rect 386 -1033 388 -993
rect 312 -1078 314 -1058
rect 479 -1063 481 -1023
rect 517 -1063 519 -1023
rect 443 -1108 445 -1088
rect 348 -1177 350 -1137
rect 386 -1177 388 -1137
rect 312 -1222 314 -1202
rect 148 -1300 150 -1260
rect 186 -1300 188 -1260
rect 6 -1393 46 -1391
rect 148 -1420 150 -1380
rect 357 -1420 359 -1380
rect 395 -1420 397 -1380
rect 511 -1380 513 -1340
rect 549 -1380 551 -1340
rect 6 -1444 46 -1442
rect 475 -1425 477 -1405
rect 321 -1465 323 -1445
rect 860 -1476 862 -1436
rect 898 -1476 900 -1436
rect 824 -1521 826 -1501
rect 357 -1564 359 -1524
rect 395 -1564 397 -1524
rect 321 -1609 323 -1589
rect 486 -1594 488 -1554
rect 524 -1594 526 -1554
rect 450 -1639 452 -1619
rect 620 -1655 622 -1615
rect 658 -1655 660 -1615
rect 360 -1734 362 -1694
rect 398 -1734 400 -1694
rect 584 -1700 586 -1680
rect 324 -1779 326 -1759
rect 491 -1764 493 -1724
rect 529 -1764 531 -1724
rect 455 -1809 457 -1789
rect 360 -1878 362 -1838
rect 398 -1878 400 -1838
rect 749 -1844 751 -1804
rect 787 -1844 789 -1804
rect 713 -1889 715 -1869
rect 324 -1923 326 -1903
rect 360 -2005 362 -1965
rect 398 -2005 400 -1965
rect 324 -2050 326 -2030
rect 491 -2035 493 -1995
rect 529 -2035 531 -1995
rect 455 -2080 457 -2060
rect 626 -2065 628 -2025
rect 664 -2065 666 -2025
rect 360 -2149 362 -2109
rect 398 -2149 400 -2109
rect 590 -2110 592 -2090
rect 324 -2194 326 -2174
<< ndiffusion >>
rect 328 262 348 263
rect 328 259 348 260
rect 377 252 378 272
rect 380 252 381 272
rect 377 220 378 240
rect 380 220 381 240
rect 328 211 348 212
rect 328 208 348 209
rect 409 193 410 213
rect 412 193 413 213
rect 115 101 116 121
rect 118 101 119 121
rect 115 69 116 89
rect 118 69 119 89
rect 382 106 383 126
rect 385 106 386 126
rect 147 68 148 88
rect 150 68 151 88
rect 185 68 186 88
rect 188 68 189 88
rect 418 76 419 96
rect 421 76 422 96
rect 456 76 457 96
rect 459 76 460 96
rect 564 81 584 82
rect 564 78 584 79
rect 613 71 614 91
rect 616 71 617 91
rect 613 39 614 59
rect 616 39 617 59
rect 564 30 584 31
rect 66 17 86 18
rect 66 14 86 15
rect 115 7 116 27
rect 118 7 119 27
rect 115 -25 116 -5
rect 118 -25 119 -5
rect 276 -22 277 -2
rect 279 -22 280 -2
rect 564 27 584 28
rect 645 12 646 32
rect 648 12 649 32
rect 66 -34 86 -33
rect 66 -37 86 -36
rect 147 -52 148 -32
rect 150 -52 151 -32
rect 312 -52 313 -32
rect 315 -52 316 -32
rect 350 -52 351 -32
rect 353 -52 354 -32
rect 115 -189 116 -169
rect 118 -189 119 -169
rect 115 -221 116 -201
rect 118 -221 119 -201
rect 459 -184 460 -164
rect 462 -184 463 -164
rect 147 -222 148 -202
rect 150 -222 151 -202
rect 185 -222 186 -202
rect 188 -222 189 -202
rect 495 -214 496 -194
rect 498 -214 499 -194
rect 533 -214 534 -194
rect 536 -214 537 -194
rect 66 -273 86 -272
rect 66 -276 86 -275
rect 115 -283 116 -263
rect 118 -283 119 -263
rect 115 -315 116 -295
rect 118 -315 119 -295
rect 356 -312 357 -292
rect 359 -312 360 -292
rect 66 -324 86 -323
rect 66 -327 86 -326
rect 147 -342 148 -322
rect 150 -342 151 -322
rect 579 -306 580 -286
rect 582 -306 583 -286
rect 392 -342 393 -322
rect 395 -342 396 -322
rect 430 -342 431 -322
rect 433 -342 434 -322
rect 615 -336 616 -316
rect 618 -336 619 -316
rect 653 -336 654 -316
rect 656 -336 657 -316
rect 766 -331 786 -330
rect 766 -334 786 -333
rect 815 -341 816 -321
rect 818 -341 819 -321
rect 815 -373 816 -353
rect 818 -373 819 -353
rect 766 -382 786 -381
rect 284 -438 285 -418
rect 287 -438 288 -418
rect 766 -385 786 -384
rect 847 -400 848 -380
rect 850 -400 851 -380
rect 320 -468 321 -448
rect 323 -468 324 -448
rect 358 -468 359 -448
rect 361 -468 362 -448
rect 413 -468 414 -448
rect 416 -468 417 -448
rect 449 -498 450 -478
rect 452 -498 453 -478
rect 487 -498 488 -478
rect 490 -498 491 -478
rect 115 -606 116 -586
rect 118 -606 119 -586
rect 115 -638 116 -618
rect 118 -638 119 -618
rect 616 -601 617 -581
rect 619 -601 620 -581
rect 147 -639 148 -619
rect 150 -639 151 -619
rect 185 -639 186 -619
rect 188 -639 189 -619
rect 652 -631 653 -611
rect 655 -631 656 -611
rect 690 -631 691 -611
rect 693 -631 694 -611
rect 66 -690 86 -689
rect 66 -693 86 -692
rect 115 -700 116 -680
rect 118 -700 119 -680
rect 115 -732 116 -712
rect 118 -732 119 -712
rect 308 -729 309 -709
rect 311 -729 312 -709
rect 66 -741 86 -740
rect 66 -744 86 -743
rect 147 -759 148 -739
rect 150 -759 151 -739
rect 783 -738 784 -718
rect 786 -738 787 -718
rect 344 -759 345 -739
rect 347 -759 348 -739
rect 382 -759 383 -739
rect 385 -759 386 -739
rect 819 -768 820 -748
rect 822 -768 823 -748
rect 857 -768 858 -748
rect 860 -768 861 -748
rect 965 -763 985 -762
rect 965 -766 985 -765
rect 1014 -773 1015 -753
rect 1017 -773 1018 -753
rect 1014 -805 1015 -785
rect 1017 -805 1018 -785
rect 965 -814 985 -813
rect 965 -817 985 -816
rect 308 -873 309 -853
rect 311 -873 312 -853
rect 1046 -832 1047 -812
rect 1049 -832 1050 -812
rect 344 -903 345 -883
rect 347 -903 348 -883
rect 382 -903 383 -883
rect 385 -903 386 -883
rect 437 -903 438 -883
rect 440 -903 441 -883
rect 473 -933 474 -913
rect 476 -933 477 -913
rect 511 -933 512 -913
rect 514 -933 515 -913
rect 612 -957 613 -937
rect 615 -957 616 -937
rect 648 -987 649 -967
rect 651 -987 652 -967
rect 686 -987 687 -967
rect 689 -987 690 -967
rect 311 -1043 312 -1023
rect 314 -1043 315 -1023
rect 347 -1073 348 -1053
rect 350 -1073 351 -1053
rect 385 -1073 386 -1053
rect 388 -1073 389 -1053
rect 442 -1073 443 -1053
rect 445 -1073 446 -1053
rect 478 -1103 479 -1083
rect 481 -1103 482 -1083
rect 516 -1103 517 -1083
rect 519 -1103 520 -1083
rect 311 -1187 312 -1167
rect 314 -1187 315 -1167
rect 347 -1217 348 -1197
rect 350 -1217 351 -1197
rect 385 -1217 386 -1197
rect 388 -1217 389 -1197
rect 115 -1307 116 -1287
rect 118 -1307 119 -1287
rect 115 -1339 116 -1319
rect 118 -1339 119 -1319
rect 147 -1340 148 -1320
rect 150 -1340 151 -1320
rect 185 -1340 186 -1320
rect 188 -1340 189 -1320
rect 66 -1391 86 -1390
rect 66 -1394 86 -1393
rect 115 -1401 116 -1381
rect 118 -1401 119 -1381
rect 115 -1433 116 -1413
rect 118 -1433 119 -1413
rect 320 -1430 321 -1410
rect 323 -1430 324 -1410
rect 474 -1390 475 -1370
rect 477 -1390 478 -1370
rect 66 -1442 86 -1441
rect 66 -1445 86 -1444
rect 147 -1460 148 -1440
rect 150 -1460 151 -1440
rect 510 -1420 511 -1400
rect 513 -1420 514 -1400
rect 548 -1420 549 -1400
rect 551 -1420 552 -1400
rect 356 -1460 357 -1440
rect 359 -1460 360 -1440
rect 394 -1460 395 -1440
rect 397 -1460 398 -1440
rect 823 -1486 824 -1466
rect 826 -1486 827 -1466
rect 859 -1516 860 -1496
rect 862 -1516 863 -1496
rect 897 -1516 898 -1496
rect 900 -1516 901 -1496
rect 320 -1574 321 -1554
rect 323 -1574 324 -1554
rect 356 -1604 357 -1584
rect 359 -1604 360 -1584
rect 394 -1604 395 -1584
rect 397 -1604 398 -1584
rect 449 -1604 450 -1584
rect 452 -1604 453 -1584
rect 485 -1634 486 -1614
rect 488 -1634 489 -1614
rect 523 -1634 524 -1614
rect 526 -1634 527 -1614
rect 583 -1665 584 -1645
rect 586 -1665 587 -1645
rect 323 -1744 324 -1724
rect 326 -1744 327 -1724
rect 619 -1695 620 -1675
rect 622 -1695 623 -1675
rect 657 -1695 658 -1675
rect 660 -1695 661 -1675
rect 359 -1774 360 -1754
rect 362 -1774 363 -1754
rect 397 -1774 398 -1754
rect 400 -1774 401 -1754
rect 454 -1774 455 -1754
rect 457 -1774 458 -1754
rect 490 -1804 491 -1784
rect 493 -1804 494 -1784
rect 528 -1804 529 -1784
rect 531 -1804 532 -1784
rect 323 -1888 324 -1868
rect 326 -1888 327 -1868
rect 712 -1854 713 -1834
rect 715 -1854 716 -1834
rect 748 -1884 749 -1864
rect 751 -1884 752 -1864
rect 786 -1884 787 -1864
rect 789 -1884 790 -1864
rect 359 -1918 360 -1898
rect 362 -1918 363 -1898
rect 397 -1918 398 -1898
rect 400 -1918 401 -1898
rect 323 -2015 324 -1995
rect 326 -2015 327 -1995
rect 359 -2045 360 -2025
rect 362 -2045 363 -2025
rect 397 -2045 398 -2025
rect 400 -2045 401 -2025
rect 454 -2045 455 -2025
rect 457 -2045 458 -2025
rect 490 -2075 491 -2055
rect 493 -2075 494 -2055
rect 528 -2075 529 -2055
rect 531 -2075 532 -2055
rect 589 -2075 590 -2055
rect 592 -2075 593 -2055
rect 323 -2159 324 -2139
rect 326 -2159 327 -2139
rect 625 -2105 626 -2085
rect 628 -2105 629 -2085
rect 663 -2105 664 -2085
rect 666 -2105 667 -2085
rect 359 -2189 360 -2169
rect 362 -2189 363 -2169
rect 397 -2189 398 -2169
rect 400 -2189 401 -2169
<< pdiffusion >>
rect 268 262 308 263
rect 268 259 308 260
rect 409 233 410 273
rect 412 233 413 273
rect 268 211 308 212
rect 268 208 308 209
rect 147 108 148 148
rect 150 108 151 148
rect 185 108 186 148
rect 188 108 189 148
rect 418 116 419 156
rect 421 116 422 156
rect 456 116 457 156
rect 459 116 460 156
rect 382 71 383 91
rect 385 71 386 91
rect 504 81 544 82
rect 504 78 544 79
rect 645 52 646 92
rect 648 52 649 92
rect 504 30 544 31
rect 6 17 46 18
rect 6 14 46 15
rect 147 -12 148 28
rect 150 -12 151 28
rect 6 -34 46 -33
rect 312 -12 313 28
rect 315 -12 316 28
rect 350 -12 351 28
rect 353 -12 354 28
rect 504 27 544 28
rect 6 -37 46 -36
rect 276 -57 277 -37
rect 279 -57 280 -37
rect 147 -182 148 -142
rect 150 -182 151 -142
rect 185 -182 186 -142
rect 188 -182 189 -142
rect 495 -174 496 -134
rect 498 -174 499 -134
rect 533 -174 534 -134
rect 536 -174 537 -134
rect 459 -219 460 -199
rect 462 -219 463 -199
rect 6 -273 46 -272
rect 6 -276 46 -275
rect 147 -302 148 -262
rect 150 -302 151 -262
rect 6 -324 46 -323
rect 392 -302 393 -262
rect 395 -302 396 -262
rect 430 -302 431 -262
rect 433 -302 434 -262
rect 6 -327 46 -326
rect 615 -296 616 -256
rect 618 -296 619 -256
rect 653 -296 654 -256
rect 656 -296 657 -256
rect 356 -347 357 -327
rect 359 -347 360 -327
rect 579 -341 580 -321
rect 582 -341 583 -321
rect 706 -331 746 -330
rect 706 -334 746 -333
rect 847 -360 848 -320
rect 850 -360 851 -320
rect 706 -382 746 -381
rect 706 -385 746 -384
rect 320 -428 321 -388
rect 323 -428 324 -388
rect 358 -428 359 -388
rect 361 -428 362 -388
rect 284 -473 285 -453
rect 287 -473 288 -453
rect 449 -458 450 -418
rect 452 -458 453 -418
rect 487 -458 488 -418
rect 490 -458 491 -418
rect 413 -503 414 -483
rect 416 -503 417 -483
rect 147 -599 148 -559
rect 150 -599 151 -559
rect 185 -599 186 -559
rect 188 -599 189 -559
rect 652 -591 653 -551
rect 655 -591 656 -551
rect 690 -591 691 -551
rect 693 -591 694 -551
rect 616 -636 617 -616
rect 619 -636 620 -616
rect 6 -690 46 -689
rect 6 -693 46 -692
rect 147 -719 148 -679
rect 150 -719 151 -679
rect 6 -741 46 -740
rect 344 -719 345 -679
rect 347 -719 348 -679
rect 382 -719 383 -679
rect 385 -719 386 -679
rect 6 -744 46 -743
rect 819 -728 820 -688
rect 822 -728 823 -688
rect 857 -728 858 -688
rect 860 -728 861 -688
rect 308 -764 309 -744
rect 311 -764 312 -744
rect 783 -773 784 -753
rect 786 -773 787 -753
rect 905 -763 945 -762
rect 905 -766 945 -765
rect 1046 -792 1047 -752
rect 1049 -792 1050 -752
rect 905 -814 945 -813
rect 905 -817 945 -816
rect 344 -863 345 -823
rect 347 -863 348 -823
rect 382 -863 383 -823
rect 385 -863 386 -823
rect 308 -908 309 -888
rect 311 -908 312 -888
rect 473 -893 474 -853
rect 476 -893 477 -853
rect 511 -893 512 -853
rect 514 -893 515 -853
rect 437 -938 438 -918
rect 440 -938 441 -918
rect 648 -947 649 -907
rect 651 -947 652 -907
rect 686 -947 687 -907
rect 689 -947 690 -907
rect 612 -992 613 -972
rect 615 -992 616 -972
rect 347 -1033 348 -993
rect 350 -1033 351 -993
rect 385 -1033 386 -993
rect 388 -1033 389 -993
rect 311 -1078 312 -1058
rect 314 -1078 315 -1058
rect 478 -1063 479 -1023
rect 481 -1063 482 -1023
rect 516 -1063 517 -1023
rect 519 -1063 520 -1023
rect 442 -1108 443 -1088
rect 445 -1108 446 -1088
rect 347 -1177 348 -1137
rect 350 -1177 351 -1137
rect 385 -1177 386 -1137
rect 388 -1177 389 -1137
rect 311 -1222 312 -1202
rect 314 -1222 315 -1202
rect 147 -1300 148 -1260
rect 150 -1300 151 -1260
rect 185 -1300 186 -1260
rect 188 -1300 189 -1260
rect 6 -1391 46 -1390
rect 6 -1394 46 -1393
rect 147 -1420 148 -1380
rect 150 -1420 151 -1380
rect 6 -1442 46 -1441
rect 356 -1420 357 -1380
rect 359 -1420 360 -1380
rect 394 -1420 395 -1380
rect 397 -1420 398 -1380
rect 510 -1380 511 -1340
rect 513 -1380 514 -1340
rect 548 -1380 549 -1340
rect 551 -1380 552 -1340
rect 6 -1445 46 -1444
rect 474 -1425 475 -1405
rect 477 -1425 478 -1405
rect 320 -1465 321 -1445
rect 323 -1465 324 -1445
rect 859 -1476 860 -1436
rect 862 -1476 863 -1436
rect 897 -1476 898 -1436
rect 900 -1476 901 -1436
rect 823 -1521 824 -1501
rect 826 -1521 827 -1501
rect 356 -1564 357 -1524
rect 359 -1564 360 -1524
rect 394 -1564 395 -1524
rect 397 -1564 398 -1524
rect 320 -1609 321 -1589
rect 323 -1609 324 -1589
rect 485 -1594 486 -1554
rect 488 -1594 489 -1554
rect 523 -1594 524 -1554
rect 526 -1594 527 -1554
rect 449 -1639 450 -1619
rect 452 -1639 453 -1619
rect 619 -1655 620 -1615
rect 622 -1655 623 -1615
rect 657 -1655 658 -1615
rect 660 -1655 661 -1615
rect 359 -1734 360 -1694
rect 362 -1734 363 -1694
rect 397 -1734 398 -1694
rect 400 -1734 401 -1694
rect 583 -1700 584 -1680
rect 586 -1700 587 -1680
rect 323 -1779 324 -1759
rect 326 -1779 327 -1759
rect 490 -1764 491 -1724
rect 493 -1764 494 -1724
rect 528 -1764 529 -1724
rect 531 -1764 532 -1724
rect 454 -1809 455 -1789
rect 457 -1809 458 -1789
rect 359 -1878 360 -1838
rect 362 -1878 363 -1838
rect 397 -1878 398 -1838
rect 400 -1878 401 -1838
rect 748 -1844 749 -1804
rect 751 -1844 752 -1804
rect 786 -1844 787 -1804
rect 789 -1844 790 -1804
rect 712 -1889 713 -1869
rect 715 -1889 716 -1869
rect 323 -1923 324 -1903
rect 326 -1923 327 -1903
rect 359 -2005 360 -1965
rect 362 -2005 363 -1965
rect 397 -2005 398 -1965
rect 400 -2005 401 -1965
rect 323 -2050 324 -2030
rect 326 -2050 327 -2030
rect 490 -2035 491 -1995
rect 493 -2035 494 -1995
rect 528 -2035 529 -1995
rect 531 -2035 532 -1995
rect 454 -2080 455 -2060
rect 457 -2080 458 -2060
rect 625 -2065 626 -2025
rect 628 -2065 629 -2025
rect 663 -2065 664 -2025
rect 666 -2065 667 -2025
rect 359 -2149 360 -2109
rect 362 -2149 363 -2109
rect 397 -2149 398 -2109
rect 400 -2149 401 -2109
rect 589 -2110 590 -2090
rect 592 -2110 593 -2090
rect 323 -2194 324 -2174
rect 326 -2194 327 -2174
<< ndcontact >>
rect 328 263 348 267
rect 328 255 348 259
rect 373 252 377 272
rect 381 252 385 272
rect 373 220 377 240
rect 381 220 385 240
rect 328 212 348 216
rect 328 204 348 208
rect 405 193 409 213
rect 413 193 417 213
rect 111 101 115 121
rect 119 101 123 121
rect 111 69 115 89
rect 119 69 123 89
rect 378 106 382 126
rect 386 106 390 126
rect 143 68 147 88
rect 151 68 155 88
rect 181 68 185 88
rect 189 68 193 88
rect 414 76 418 96
rect 422 76 426 96
rect 452 76 456 96
rect 460 76 464 96
rect 564 82 584 86
rect 564 74 584 78
rect 609 71 613 91
rect 617 71 621 91
rect 609 39 613 59
rect 617 39 621 59
rect 564 31 584 35
rect 66 18 86 22
rect 66 10 86 14
rect 111 7 115 27
rect 119 7 123 27
rect 111 -25 115 -5
rect 119 -25 123 -5
rect 66 -33 86 -29
rect 272 -22 276 -2
rect 280 -22 284 -2
rect 564 23 584 27
rect 641 12 645 32
rect 649 12 653 32
rect 66 -41 86 -37
rect 143 -52 147 -32
rect 151 -52 155 -32
rect 308 -52 312 -32
rect 316 -52 320 -32
rect 346 -52 350 -32
rect 354 -52 358 -32
rect 111 -189 115 -169
rect 119 -189 123 -169
rect 111 -221 115 -201
rect 119 -221 123 -201
rect 455 -184 459 -164
rect 463 -184 467 -164
rect 143 -222 147 -202
rect 151 -222 155 -202
rect 181 -222 185 -202
rect 189 -222 193 -202
rect 491 -214 495 -194
rect 499 -214 503 -194
rect 529 -214 533 -194
rect 537 -214 541 -194
rect 66 -272 86 -268
rect 66 -280 86 -276
rect 111 -283 115 -263
rect 119 -283 123 -263
rect 111 -315 115 -295
rect 119 -315 123 -295
rect 66 -323 86 -319
rect 352 -312 356 -292
rect 360 -312 364 -292
rect 66 -331 86 -327
rect 143 -342 147 -322
rect 151 -342 155 -322
rect 575 -306 579 -286
rect 583 -306 587 -286
rect 388 -342 392 -322
rect 396 -342 400 -322
rect 426 -342 430 -322
rect 434 -342 438 -322
rect 611 -336 615 -316
rect 619 -336 623 -316
rect 649 -336 653 -316
rect 657 -336 661 -316
rect 766 -330 786 -326
rect 766 -338 786 -334
rect 811 -341 815 -321
rect 819 -341 823 -321
rect 811 -373 815 -353
rect 819 -373 823 -353
rect 766 -381 786 -377
rect 280 -438 284 -418
rect 288 -438 292 -418
rect 766 -389 786 -385
rect 843 -400 847 -380
rect 851 -400 855 -380
rect 316 -468 320 -448
rect 324 -468 328 -448
rect 354 -468 358 -448
rect 362 -468 366 -448
rect 409 -468 413 -448
rect 417 -468 421 -448
rect 445 -498 449 -478
rect 453 -498 457 -478
rect 483 -498 487 -478
rect 491 -498 495 -478
rect 111 -606 115 -586
rect 119 -606 123 -586
rect 111 -638 115 -618
rect 119 -638 123 -618
rect 612 -601 616 -581
rect 620 -601 624 -581
rect 143 -639 147 -619
rect 151 -639 155 -619
rect 181 -639 185 -619
rect 189 -639 193 -619
rect 648 -631 652 -611
rect 656 -631 660 -611
rect 686 -631 690 -611
rect 694 -631 698 -611
rect 66 -689 86 -685
rect 66 -697 86 -693
rect 111 -700 115 -680
rect 119 -700 123 -680
rect 111 -732 115 -712
rect 119 -732 123 -712
rect 66 -740 86 -736
rect 304 -729 308 -709
rect 312 -729 316 -709
rect 66 -748 86 -744
rect 143 -759 147 -739
rect 151 -759 155 -739
rect 779 -738 783 -718
rect 787 -738 791 -718
rect 340 -759 344 -739
rect 348 -759 352 -739
rect 378 -759 382 -739
rect 386 -759 390 -739
rect 815 -768 819 -748
rect 823 -768 827 -748
rect 853 -768 857 -748
rect 861 -768 865 -748
rect 965 -762 985 -758
rect 965 -770 985 -766
rect 1010 -773 1014 -753
rect 1018 -773 1022 -753
rect 1010 -805 1014 -785
rect 1018 -805 1022 -785
rect 965 -813 985 -809
rect 965 -821 985 -817
rect 304 -873 308 -853
rect 312 -873 316 -853
rect 1042 -832 1046 -812
rect 1050 -832 1054 -812
rect 340 -903 344 -883
rect 348 -903 352 -883
rect 378 -903 382 -883
rect 386 -903 390 -883
rect 433 -903 437 -883
rect 441 -903 445 -883
rect 469 -933 473 -913
rect 477 -933 481 -913
rect 507 -933 511 -913
rect 515 -933 519 -913
rect 608 -957 612 -937
rect 616 -957 620 -937
rect 644 -987 648 -967
rect 652 -987 656 -967
rect 682 -987 686 -967
rect 690 -987 694 -967
rect 307 -1043 311 -1023
rect 315 -1043 319 -1023
rect 343 -1073 347 -1053
rect 351 -1073 355 -1053
rect 381 -1073 385 -1053
rect 389 -1073 393 -1053
rect 438 -1073 442 -1053
rect 446 -1073 450 -1053
rect 474 -1103 478 -1083
rect 482 -1103 486 -1083
rect 512 -1103 516 -1083
rect 520 -1103 524 -1083
rect 307 -1187 311 -1167
rect 315 -1187 319 -1167
rect 343 -1217 347 -1197
rect 351 -1217 355 -1197
rect 381 -1217 385 -1197
rect 389 -1217 393 -1197
rect 111 -1307 115 -1287
rect 119 -1307 123 -1287
rect 111 -1339 115 -1319
rect 119 -1339 123 -1319
rect 143 -1340 147 -1320
rect 151 -1340 155 -1320
rect 181 -1340 185 -1320
rect 189 -1340 193 -1320
rect 66 -1390 86 -1386
rect 66 -1398 86 -1394
rect 111 -1401 115 -1381
rect 119 -1401 123 -1381
rect 111 -1433 115 -1413
rect 119 -1433 123 -1413
rect 66 -1441 86 -1437
rect 316 -1430 320 -1410
rect 324 -1430 328 -1410
rect 470 -1390 474 -1370
rect 478 -1390 482 -1370
rect 66 -1449 86 -1445
rect 143 -1460 147 -1440
rect 151 -1460 155 -1440
rect 506 -1420 510 -1400
rect 514 -1420 518 -1400
rect 544 -1420 548 -1400
rect 552 -1420 556 -1400
rect 352 -1460 356 -1440
rect 360 -1460 364 -1440
rect 390 -1460 394 -1440
rect 398 -1460 402 -1440
rect 819 -1486 823 -1466
rect 827 -1486 831 -1466
rect 855 -1516 859 -1496
rect 863 -1516 867 -1496
rect 893 -1516 897 -1496
rect 901 -1516 905 -1496
rect 316 -1574 320 -1554
rect 324 -1574 328 -1554
rect 352 -1604 356 -1584
rect 360 -1604 364 -1584
rect 390 -1604 394 -1584
rect 398 -1604 402 -1584
rect 445 -1604 449 -1584
rect 453 -1604 457 -1584
rect 481 -1634 485 -1614
rect 489 -1634 493 -1614
rect 519 -1634 523 -1614
rect 527 -1634 531 -1614
rect 579 -1665 583 -1645
rect 587 -1665 591 -1645
rect 319 -1744 323 -1724
rect 327 -1744 331 -1724
rect 615 -1695 619 -1675
rect 623 -1695 627 -1675
rect 653 -1695 657 -1675
rect 661 -1695 665 -1675
rect 355 -1774 359 -1754
rect 363 -1774 367 -1754
rect 393 -1774 397 -1754
rect 401 -1774 405 -1754
rect 450 -1774 454 -1754
rect 458 -1774 462 -1754
rect 486 -1804 490 -1784
rect 494 -1804 498 -1784
rect 524 -1804 528 -1784
rect 532 -1804 536 -1784
rect 319 -1888 323 -1868
rect 327 -1888 331 -1868
rect 708 -1854 712 -1834
rect 716 -1854 720 -1834
rect 744 -1884 748 -1864
rect 752 -1884 756 -1864
rect 782 -1884 786 -1864
rect 790 -1884 794 -1864
rect 355 -1918 359 -1898
rect 363 -1918 367 -1898
rect 393 -1918 397 -1898
rect 401 -1918 405 -1898
rect 319 -2015 323 -1995
rect 327 -2015 331 -1995
rect 355 -2045 359 -2025
rect 363 -2045 367 -2025
rect 393 -2045 397 -2025
rect 401 -2045 405 -2025
rect 450 -2045 454 -2025
rect 458 -2045 462 -2025
rect 486 -2075 490 -2055
rect 494 -2075 498 -2055
rect 524 -2075 528 -2055
rect 532 -2075 536 -2055
rect 585 -2075 589 -2055
rect 593 -2075 597 -2055
rect 319 -2159 323 -2139
rect 327 -2159 331 -2139
rect 621 -2105 625 -2085
rect 629 -2105 633 -2085
rect 659 -2105 663 -2085
rect 667 -2105 671 -2085
rect 355 -2189 359 -2169
rect 363 -2189 367 -2169
rect 393 -2189 397 -2169
rect 401 -2189 405 -2169
<< pdcontact >>
rect 268 263 308 267
rect 268 255 308 259
rect 405 233 409 273
rect 413 233 417 273
rect 268 212 308 216
rect 268 204 308 208
rect 143 108 147 148
rect 151 108 155 148
rect 181 108 185 148
rect 189 108 193 148
rect 414 116 418 156
rect 422 116 426 156
rect 452 116 456 156
rect 460 116 464 156
rect 378 71 382 91
rect 386 71 390 91
rect 504 82 544 86
rect 504 74 544 78
rect 641 52 645 92
rect 649 52 653 92
rect 504 31 544 35
rect 6 18 46 22
rect 6 10 46 14
rect 143 -12 147 28
rect 151 -12 155 28
rect 6 -33 46 -29
rect 308 -12 312 28
rect 316 -12 320 28
rect 346 -12 350 28
rect 354 -12 358 28
rect 504 23 544 27
rect 6 -41 46 -37
rect 272 -57 276 -37
rect 280 -57 284 -37
rect 143 -182 147 -142
rect 151 -182 155 -142
rect 181 -182 185 -142
rect 189 -182 193 -142
rect 491 -174 495 -134
rect 499 -174 503 -134
rect 529 -174 533 -134
rect 537 -174 541 -134
rect 455 -219 459 -199
rect 463 -219 467 -199
rect 6 -272 46 -268
rect 6 -280 46 -276
rect 143 -302 147 -262
rect 151 -302 155 -262
rect 6 -323 46 -319
rect 388 -302 392 -262
rect 396 -302 400 -262
rect 426 -302 430 -262
rect 434 -302 438 -262
rect 6 -331 46 -327
rect 611 -296 615 -256
rect 619 -296 623 -256
rect 649 -296 653 -256
rect 657 -296 661 -256
rect 352 -347 356 -327
rect 360 -347 364 -327
rect 575 -341 579 -321
rect 583 -341 587 -321
rect 706 -330 746 -326
rect 706 -338 746 -334
rect 843 -360 847 -320
rect 851 -360 855 -320
rect 706 -381 746 -377
rect 316 -428 320 -388
rect 324 -428 328 -388
rect 354 -428 358 -388
rect 362 -428 366 -388
rect 706 -389 746 -385
rect 280 -473 284 -453
rect 288 -473 292 -453
rect 445 -458 449 -418
rect 453 -458 457 -418
rect 483 -458 487 -418
rect 491 -458 495 -418
rect 409 -503 413 -483
rect 417 -503 421 -483
rect 143 -599 147 -559
rect 151 -599 155 -559
rect 181 -599 185 -559
rect 189 -599 193 -559
rect 648 -591 652 -551
rect 656 -591 660 -551
rect 686 -591 690 -551
rect 694 -591 698 -551
rect 612 -636 616 -616
rect 620 -636 624 -616
rect 6 -689 46 -685
rect 6 -697 46 -693
rect 143 -719 147 -679
rect 151 -719 155 -679
rect 6 -740 46 -736
rect 340 -719 344 -679
rect 348 -719 352 -679
rect 378 -719 382 -679
rect 386 -719 390 -679
rect 6 -748 46 -744
rect 815 -728 819 -688
rect 823 -728 827 -688
rect 853 -728 857 -688
rect 861 -728 865 -688
rect 304 -764 308 -744
rect 312 -764 316 -744
rect 779 -773 783 -753
rect 787 -773 791 -753
rect 905 -762 945 -758
rect 905 -770 945 -766
rect 1042 -792 1046 -752
rect 1050 -792 1054 -752
rect 905 -813 945 -809
rect 905 -821 945 -817
rect 340 -863 344 -823
rect 348 -863 352 -823
rect 378 -863 382 -823
rect 386 -863 390 -823
rect 304 -908 308 -888
rect 312 -908 316 -888
rect 469 -893 473 -853
rect 477 -893 481 -853
rect 507 -893 511 -853
rect 515 -893 519 -853
rect 433 -938 437 -918
rect 441 -938 445 -918
rect 644 -947 648 -907
rect 652 -947 656 -907
rect 682 -947 686 -907
rect 690 -947 694 -907
rect 608 -992 612 -972
rect 616 -992 620 -972
rect 343 -1033 347 -993
rect 351 -1033 355 -993
rect 381 -1033 385 -993
rect 389 -1033 393 -993
rect 307 -1078 311 -1058
rect 315 -1078 319 -1058
rect 474 -1063 478 -1023
rect 482 -1063 486 -1023
rect 512 -1063 516 -1023
rect 520 -1063 524 -1023
rect 438 -1108 442 -1088
rect 446 -1108 450 -1088
rect 343 -1177 347 -1137
rect 351 -1177 355 -1137
rect 381 -1177 385 -1137
rect 389 -1177 393 -1137
rect 307 -1222 311 -1202
rect 315 -1222 319 -1202
rect 143 -1300 147 -1260
rect 151 -1300 155 -1260
rect 181 -1300 185 -1260
rect 189 -1300 193 -1260
rect 6 -1390 46 -1386
rect 6 -1398 46 -1394
rect 143 -1420 147 -1380
rect 151 -1420 155 -1380
rect 6 -1441 46 -1437
rect 352 -1420 356 -1380
rect 360 -1420 364 -1380
rect 390 -1420 394 -1380
rect 398 -1420 402 -1380
rect 506 -1380 510 -1340
rect 514 -1380 518 -1340
rect 544 -1380 548 -1340
rect 552 -1380 556 -1340
rect 6 -1449 46 -1445
rect 470 -1425 474 -1405
rect 478 -1425 482 -1405
rect 316 -1465 320 -1445
rect 324 -1465 328 -1445
rect 855 -1476 859 -1436
rect 863 -1476 867 -1436
rect 893 -1476 897 -1436
rect 901 -1476 905 -1436
rect 819 -1521 823 -1501
rect 827 -1521 831 -1501
rect 352 -1564 356 -1524
rect 360 -1564 364 -1524
rect 390 -1564 394 -1524
rect 398 -1564 402 -1524
rect 316 -1609 320 -1589
rect 324 -1609 328 -1589
rect 481 -1594 485 -1554
rect 489 -1594 493 -1554
rect 519 -1594 523 -1554
rect 527 -1594 531 -1554
rect 445 -1639 449 -1619
rect 453 -1639 457 -1619
rect 615 -1655 619 -1615
rect 623 -1655 627 -1615
rect 653 -1655 657 -1615
rect 661 -1655 665 -1615
rect 355 -1734 359 -1694
rect 363 -1734 367 -1694
rect 393 -1734 397 -1694
rect 401 -1734 405 -1694
rect 579 -1700 583 -1680
rect 587 -1700 591 -1680
rect 319 -1779 323 -1759
rect 327 -1779 331 -1759
rect 486 -1764 490 -1724
rect 494 -1764 498 -1724
rect 524 -1764 528 -1724
rect 532 -1764 536 -1724
rect 450 -1809 454 -1789
rect 458 -1809 462 -1789
rect 355 -1878 359 -1838
rect 363 -1878 367 -1838
rect 393 -1878 397 -1838
rect 401 -1878 405 -1838
rect 744 -1844 748 -1804
rect 752 -1844 756 -1804
rect 782 -1844 786 -1804
rect 790 -1844 794 -1804
rect 708 -1889 712 -1869
rect 716 -1889 720 -1869
rect 319 -1923 323 -1903
rect 327 -1923 331 -1903
rect 355 -2005 359 -1965
rect 363 -2005 367 -1965
rect 393 -2005 397 -1965
rect 401 -2005 405 -1965
rect 319 -2050 323 -2030
rect 327 -2050 331 -2030
rect 486 -2035 490 -1995
rect 494 -2035 498 -1995
rect 524 -2035 528 -1995
rect 532 -2035 536 -1995
rect 450 -2080 454 -2060
rect 458 -2080 462 -2060
rect 621 -2065 625 -2025
rect 629 -2065 633 -2025
rect 659 -2065 663 -2025
rect 667 -2065 671 -2025
rect 355 -2149 359 -2109
rect 363 -2149 367 -2109
rect 393 -2149 397 -2109
rect 401 -2149 405 -2109
rect 585 -2110 589 -2090
rect 593 -2110 597 -2090
rect 319 -2194 323 -2174
rect 327 -2194 331 -2174
<< psubstratepcontact >>
rect 357 271 361 275
rect 357 247 361 251
rect 357 220 361 224
rect 357 196 361 200
rect 397 180 401 184
rect 421 180 425 184
rect 103 62 107 66
rect 593 90 597 94
rect 593 66 597 70
rect 135 55 139 59
rect 159 55 163 59
rect 173 55 177 59
rect 197 55 201 59
rect 406 56 410 60
rect 468 56 472 60
rect 95 26 99 30
rect 593 39 597 43
rect 95 2 99 6
rect 95 -25 99 -21
rect 593 15 597 19
rect 633 -1 637 3
rect 657 -1 661 3
rect 95 -49 99 -45
rect 135 -65 139 -61
rect 159 -65 163 -61
rect 264 -72 268 -68
rect 362 -72 366 -68
rect 103 -228 107 -224
rect 135 -235 139 -231
rect 159 -235 163 -231
rect 173 -235 177 -231
rect 197 -235 201 -231
rect 483 -234 487 -230
rect 545 -234 549 -230
rect 95 -264 99 -260
rect 95 -288 99 -284
rect 95 -315 99 -311
rect 95 -339 99 -335
rect 795 -322 799 -318
rect 135 -355 139 -351
rect 159 -355 163 -351
rect 795 -346 799 -342
rect 603 -356 607 -352
rect 665 -356 669 -352
rect 344 -362 348 -358
rect 442 -362 446 -358
rect 795 -373 799 -369
rect 795 -397 799 -393
rect 835 -413 839 -409
rect 859 -413 863 -409
rect 272 -488 276 -484
rect 370 -488 374 -484
rect 401 -518 405 -514
rect 499 -518 503 -514
rect 103 -645 107 -641
rect 135 -652 139 -648
rect 159 -652 163 -648
rect 173 -652 177 -648
rect 197 -652 201 -648
rect 640 -651 644 -647
rect 702 -651 706 -647
rect 95 -681 99 -677
rect 95 -705 99 -701
rect 95 -732 99 -728
rect 95 -756 99 -752
rect 135 -772 139 -768
rect 159 -772 163 -768
rect 994 -754 998 -750
rect 296 -779 300 -775
rect 394 -779 398 -775
rect 994 -778 998 -774
rect 807 -788 811 -784
rect 869 -788 873 -784
rect 994 -805 998 -801
rect 994 -829 998 -825
rect 1034 -845 1038 -841
rect 1058 -845 1062 -841
rect 296 -923 300 -919
rect 394 -923 398 -919
rect 425 -953 429 -949
rect 523 -953 527 -949
rect 636 -1007 640 -1003
rect 698 -1007 702 -1003
rect 299 -1093 303 -1089
rect 397 -1093 401 -1089
rect 430 -1123 434 -1119
rect 528 -1123 532 -1119
rect 299 -1237 303 -1233
rect 397 -1237 401 -1233
rect 103 -1346 107 -1342
rect 135 -1353 139 -1349
rect 159 -1353 163 -1349
rect 173 -1353 177 -1349
rect 197 -1353 201 -1349
rect 95 -1382 99 -1378
rect 95 -1406 99 -1402
rect 95 -1433 99 -1429
rect 95 -1457 99 -1453
rect 498 -1440 502 -1436
rect 560 -1440 564 -1436
rect 135 -1473 139 -1469
rect 159 -1473 163 -1469
rect 308 -1480 312 -1476
rect 406 -1480 410 -1476
rect 847 -1536 851 -1532
rect 909 -1536 913 -1532
rect 308 -1624 312 -1620
rect 406 -1624 410 -1620
rect 437 -1654 441 -1650
rect 535 -1654 539 -1650
rect 607 -1715 611 -1711
rect 669 -1715 673 -1711
rect 311 -1794 315 -1790
rect 409 -1794 413 -1790
rect 442 -1824 446 -1820
rect 540 -1824 544 -1820
rect 736 -1904 740 -1900
rect 798 -1904 802 -1900
rect 311 -1938 315 -1934
rect 409 -1938 413 -1934
rect 311 -2065 315 -2061
rect 409 -2065 413 -2061
rect 442 -2095 446 -2091
rect 540 -2095 544 -2091
rect 577 -2125 581 -2121
rect 675 -2125 679 -2121
rect 311 -2209 315 -2205
rect 409 -2209 413 -2205
<< nsubstratencontact >>
rect 256 270 260 274
rect 398 281 402 285
rect 420 281 424 285
rect 256 248 260 252
rect 256 219 260 223
rect 256 197 260 201
rect 407 164 411 168
rect 467 164 471 168
rect 136 156 140 160
rect 158 156 162 160
rect 174 156 178 160
rect 196 156 200 160
rect 492 89 496 93
rect 634 100 638 104
rect 656 100 660 104
rect 492 67 496 71
rect -6 25 -2 29
rect 136 36 140 40
rect 158 36 162 40
rect 301 36 305 40
rect 361 36 365 40
rect 492 38 496 42
rect -6 3 -2 7
rect -6 -26 -2 -22
rect 492 16 496 20
rect -6 -48 -2 -44
rect 484 -126 488 -122
rect 544 -126 548 -122
rect 136 -134 140 -130
rect 158 -134 162 -130
rect 174 -134 178 -130
rect 196 -134 200 -130
rect 604 -248 608 -244
rect 664 -248 668 -244
rect -6 -265 -2 -261
rect 136 -254 140 -250
rect 158 -254 162 -250
rect 381 -254 385 -250
rect 441 -254 445 -250
rect -6 -287 -2 -283
rect -6 -316 -2 -312
rect -6 -338 -2 -334
rect 694 -323 698 -319
rect 836 -312 840 -308
rect 858 -312 862 -308
rect 694 -345 698 -341
rect 694 -374 698 -370
rect 309 -380 313 -376
rect 369 -380 373 -376
rect 694 -396 698 -392
rect 438 -410 442 -406
rect 498 -410 502 -406
rect 641 -543 645 -539
rect 701 -543 705 -539
rect 136 -551 140 -547
rect 158 -551 162 -547
rect 174 -551 178 -547
rect 196 -551 200 -547
rect -6 -682 -2 -678
rect 136 -671 140 -667
rect 158 -671 162 -667
rect 333 -671 337 -667
rect 393 -671 397 -667
rect -6 -704 -2 -700
rect -6 -733 -2 -729
rect 808 -680 812 -676
rect 868 -680 872 -676
rect -6 -755 -2 -751
rect 893 -755 897 -751
rect 1035 -744 1039 -740
rect 1057 -744 1061 -740
rect 893 -777 897 -773
rect 893 -806 897 -802
rect 333 -815 337 -811
rect 393 -815 397 -811
rect 893 -828 897 -824
rect 462 -845 466 -841
rect 522 -845 526 -841
rect 637 -899 641 -895
rect 697 -899 701 -895
rect 336 -985 340 -981
rect 396 -985 400 -981
rect 467 -1015 471 -1011
rect 527 -1015 531 -1011
rect 336 -1129 340 -1125
rect 396 -1129 400 -1125
rect 136 -1252 140 -1248
rect 158 -1252 162 -1248
rect 174 -1252 178 -1248
rect 196 -1252 200 -1248
rect 499 -1332 503 -1328
rect 559 -1332 563 -1328
rect -6 -1383 -2 -1379
rect 136 -1372 140 -1368
rect 158 -1372 162 -1368
rect 345 -1372 349 -1368
rect 405 -1372 409 -1368
rect -6 -1405 -2 -1401
rect -6 -1434 -2 -1430
rect -6 -1456 -2 -1452
rect 848 -1428 852 -1424
rect 908 -1428 912 -1424
rect 345 -1516 349 -1512
rect 405 -1516 409 -1512
rect 474 -1546 478 -1542
rect 534 -1546 538 -1542
rect 608 -1607 612 -1603
rect 668 -1607 672 -1603
rect 348 -1686 352 -1682
rect 408 -1686 412 -1682
rect 479 -1716 483 -1712
rect 539 -1716 543 -1712
rect 737 -1796 741 -1792
rect 797 -1796 801 -1792
rect 348 -1830 352 -1826
rect 408 -1830 412 -1826
rect 348 -1957 352 -1953
rect 408 -1957 412 -1953
rect 479 -1987 483 -1983
rect 539 -1987 543 -1983
rect 614 -2017 618 -2013
rect 674 -2017 678 -2013
rect 348 -2101 352 -2097
rect 408 -2101 412 -2097
<< polysilicon >>
rect 378 272 380 285
rect 410 273 412 277
rect 264 260 268 262
rect 308 260 328 262
rect 348 260 352 262
rect 378 248 380 252
rect 350 242 380 244
rect 350 239 352 242
rect 378 240 380 242
rect 378 216 380 220
rect 410 213 412 233
rect 264 209 268 211
rect 308 209 328 211
rect 348 209 352 211
rect 410 189 412 193
rect 419 156 421 160
rect 457 156 459 160
rect 148 148 150 152
rect 186 148 188 152
rect 74 123 118 125
rect 116 121 118 123
rect 383 126 385 130
rect 116 97 118 101
rect 116 89 118 93
rect 148 88 150 108
rect 186 88 188 108
rect 383 91 385 106
rect 419 96 421 116
rect 457 96 459 116
rect 116 53 118 69
rect 614 91 616 104
rect 646 92 648 96
rect 500 79 504 81
rect 544 79 564 81
rect 584 79 588 81
rect 419 72 421 76
rect 457 72 459 76
rect 148 64 150 68
rect 186 64 188 68
rect 383 59 385 71
rect 614 67 616 71
rect 586 61 616 63
rect 586 58 588 61
rect 614 59 616 61
rect 49 51 118 53
rect 116 27 118 40
rect 614 35 616 39
rect 148 28 150 32
rect 313 28 315 32
rect 351 28 353 32
rect 646 32 648 52
rect 500 28 504 30
rect 544 28 564 30
rect 584 28 588 30
rect 2 15 6 17
rect 46 15 66 17
rect 86 15 90 17
rect 116 3 118 7
rect 88 -3 118 -1
rect 88 -6 90 -3
rect 116 -5 118 -3
rect 277 -2 279 6
rect 116 -29 118 -25
rect 148 -32 150 -12
rect 646 8 648 12
rect 2 -36 6 -34
rect 46 -36 66 -34
rect 86 -36 90 -34
rect 277 -37 279 -22
rect 313 -32 315 -12
rect 351 -32 353 -12
rect 148 -56 150 -52
rect 313 -56 315 -52
rect 351 -56 353 -52
rect 277 -61 279 -57
rect 496 -134 498 -130
rect 534 -134 536 -130
rect 148 -142 150 -138
rect 186 -142 188 -138
rect 74 -167 118 -165
rect 116 -169 118 -167
rect 460 -164 462 -160
rect 116 -193 118 -189
rect 116 -201 118 -197
rect 148 -202 150 -182
rect 186 -202 188 -182
rect 460 -199 462 -184
rect 496 -194 498 -174
rect 534 -194 536 -174
rect 116 -237 118 -221
rect 496 -218 498 -214
rect 534 -218 536 -214
rect 148 -226 150 -222
rect 186 -226 188 -222
rect 460 -231 462 -219
rect 49 -239 118 -237
rect 116 -263 118 -250
rect 616 -256 618 -252
rect 654 -256 656 -252
rect 148 -262 150 -258
rect 393 -262 395 -258
rect 431 -262 433 -258
rect 2 -275 6 -273
rect 46 -275 66 -273
rect 86 -275 90 -273
rect 116 -287 118 -283
rect 88 -293 118 -291
rect 88 -296 90 -293
rect 116 -295 118 -293
rect 357 -292 359 -284
rect 116 -319 118 -315
rect 148 -322 150 -302
rect 580 -286 582 -282
rect 2 -326 6 -324
rect 46 -326 66 -324
rect 86 -326 90 -324
rect 357 -327 359 -312
rect 393 -322 395 -302
rect 431 -322 433 -302
rect 580 -321 582 -306
rect 616 -316 618 -296
rect 654 -316 656 -296
rect 148 -346 150 -342
rect 816 -321 818 -308
rect 848 -320 850 -316
rect 702 -333 706 -331
rect 746 -333 766 -331
rect 786 -333 790 -331
rect 616 -340 618 -336
rect 654 -340 656 -336
rect 393 -346 395 -342
rect 431 -346 433 -342
rect 357 -351 359 -347
rect 580 -353 582 -341
rect 816 -345 818 -341
rect 788 -351 818 -349
rect 788 -354 790 -351
rect 816 -353 818 -351
rect 816 -377 818 -373
rect 848 -380 850 -360
rect 702 -384 706 -382
rect 746 -384 766 -382
rect 786 -384 790 -382
rect 321 -388 323 -384
rect 359 -388 361 -384
rect 285 -418 287 -410
rect 848 -404 850 -400
rect 450 -418 452 -414
rect 488 -418 490 -414
rect 285 -453 287 -438
rect 321 -448 323 -428
rect 359 -448 361 -428
rect 414 -448 416 -440
rect 321 -472 323 -468
rect 359 -472 361 -468
rect 285 -477 287 -473
rect 414 -483 416 -468
rect 450 -478 452 -458
rect 488 -478 490 -458
rect 450 -502 452 -498
rect 488 -502 490 -498
rect 414 -507 416 -503
rect 653 -551 655 -547
rect 691 -551 693 -547
rect 148 -559 150 -555
rect 186 -559 188 -555
rect 74 -584 118 -582
rect 116 -586 118 -584
rect 617 -581 619 -577
rect 116 -610 118 -606
rect 116 -618 118 -614
rect 148 -619 150 -599
rect 186 -619 188 -599
rect 617 -616 619 -601
rect 653 -611 655 -591
rect 691 -611 693 -591
rect 116 -654 118 -638
rect 653 -635 655 -631
rect 691 -635 693 -631
rect 148 -643 150 -639
rect 186 -643 188 -639
rect 617 -648 619 -636
rect 49 -656 118 -654
rect 116 -680 118 -667
rect 148 -679 150 -675
rect 345 -679 347 -675
rect 383 -679 385 -675
rect 2 -692 6 -690
rect 46 -692 66 -690
rect 86 -692 90 -690
rect 116 -704 118 -700
rect 88 -710 118 -708
rect 88 -713 90 -710
rect 116 -712 118 -710
rect 309 -709 311 -701
rect 116 -736 118 -732
rect 148 -739 150 -719
rect 820 -688 822 -684
rect 858 -688 860 -684
rect 784 -718 786 -714
rect 2 -743 6 -741
rect 46 -743 66 -741
rect 86 -743 90 -741
rect 309 -744 311 -729
rect 345 -739 347 -719
rect 383 -739 385 -719
rect 148 -763 150 -759
rect 784 -753 786 -738
rect 820 -748 822 -728
rect 858 -748 860 -728
rect 345 -763 347 -759
rect 383 -763 385 -759
rect 309 -768 311 -764
rect 1015 -753 1017 -740
rect 1047 -752 1049 -748
rect 901 -765 905 -763
rect 945 -765 965 -763
rect 985 -765 989 -763
rect 820 -772 822 -768
rect 858 -772 860 -768
rect 784 -785 786 -773
rect 1015 -777 1017 -773
rect 987 -783 1017 -781
rect 987 -786 989 -783
rect 1015 -785 1017 -783
rect 1015 -809 1017 -805
rect 1047 -812 1049 -792
rect 901 -816 905 -814
rect 945 -816 965 -814
rect 985 -816 989 -814
rect 345 -823 347 -819
rect 383 -823 385 -819
rect 309 -853 311 -845
rect 1047 -836 1049 -832
rect 474 -853 476 -849
rect 512 -853 514 -849
rect 309 -888 311 -873
rect 345 -883 347 -863
rect 383 -883 385 -863
rect 438 -883 440 -875
rect 345 -907 347 -903
rect 383 -907 385 -903
rect 309 -912 311 -908
rect 438 -918 440 -903
rect 474 -913 476 -893
rect 512 -913 514 -893
rect 649 -907 651 -903
rect 687 -907 689 -903
rect 474 -937 476 -933
rect 512 -937 514 -933
rect 613 -937 615 -933
rect 438 -942 440 -938
rect 613 -972 615 -957
rect 649 -967 651 -947
rect 687 -967 689 -947
rect 348 -993 350 -989
rect 386 -993 388 -989
rect 649 -991 651 -987
rect 687 -991 689 -987
rect 312 -1023 314 -1015
rect 613 -1004 615 -992
rect 479 -1023 481 -1019
rect 517 -1023 519 -1019
rect 312 -1058 314 -1043
rect 348 -1053 350 -1033
rect 386 -1053 388 -1033
rect 443 -1053 445 -1045
rect 348 -1077 350 -1073
rect 386 -1077 388 -1073
rect 312 -1082 314 -1078
rect 443 -1088 445 -1073
rect 479 -1083 481 -1063
rect 517 -1083 519 -1063
rect 479 -1107 481 -1103
rect 517 -1107 519 -1103
rect 443 -1112 445 -1108
rect 348 -1137 350 -1133
rect 386 -1137 388 -1133
rect 312 -1167 314 -1159
rect 312 -1202 314 -1187
rect 348 -1197 350 -1177
rect 386 -1197 388 -1177
rect 348 -1221 350 -1217
rect 386 -1221 388 -1217
rect 312 -1226 314 -1222
rect 148 -1260 150 -1256
rect 186 -1260 188 -1256
rect 74 -1285 118 -1283
rect 116 -1287 118 -1285
rect 116 -1311 118 -1307
rect 116 -1319 118 -1315
rect 148 -1320 150 -1300
rect 186 -1320 188 -1300
rect 116 -1355 118 -1339
rect 511 -1340 513 -1336
rect 549 -1340 551 -1336
rect 148 -1344 150 -1340
rect 186 -1344 188 -1340
rect 49 -1357 118 -1355
rect 116 -1381 118 -1368
rect 475 -1370 477 -1366
rect 148 -1380 150 -1376
rect 357 -1380 359 -1376
rect 395 -1380 397 -1376
rect 2 -1393 6 -1391
rect 46 -1393 66 -1391
rect 86 -1393 90 -1391
rect 116 -1405 118 -1401
rect 88 -1411 118 -1409
rect 88 -1414 90 -1411
rect 116 -1413 118 -1411
rect 321 -1410 323 -1402
rect 116 -1437 118 -1433
rect 148 -1440 150 -1420
rect 475 -1405 477 -1390
rect 511 -1400 513 -1380
rect 549 -1400 551 -1380
rect 2 -1444 6 -1442
rect 46 -1444 66 -1442
rect 86 -1444 90 -1442
rect 321 -1445 323 -1430
rect 357 -1440 359 -1420
rect 395 -1440 397 -1420
rect 511 -1424 513 -1420
rect 549 -1424 551 -1420
rect 475 -1437 477 -1425
rect 860 -1436 862 -1432
rect 898 -1436 900 -1432
rect 148 -1464 150 -1460
rect 357 -1464 359 -1460
rect 395 -1464 397 -1460
rect 321 -1469 323 -1465
rect 824 -1466 826 -1462
rect 824 -1501 826 -1486
rect 860 -1496 862 -1476
rect 898 -1496 900 -1476
rect 357 -1524 359 -1520
rect 395 -1524 397 -1520
rect 860 -1520 862 -1516
rect 898 -1520 900 -1516
rect 321 -1554 323 -1546
rect 824 -1533 826 -1521
rect 486 -1554 488 -1550
rect 524 -1554 526 -1550
rect 321 -1589 323 -1574
rect 357 -1584 359 -1564
rect 395 -1584 397 -1564
rect 450 -1584 452 -1576
rect 357 -1608 359 -1604
rect 395 -1608 397 -1604
rect 321 -1613 323 -1609
rect 450 -1619 452 -1604
rect 486 -1614 488 -1594
rect 524 -1614 526 -1594
rect 620 -1615 622 -1611
rect 658 -1615 660 -1611
rect 486 -1638 488 -1634
rect 524 -1638 526 -1634
rect 450 -1643 452 -1639
rect 584 -1645 586 -1641
rect 584 -1680 586 -1665
rect 620 -1675 622 -1655
rect 658 -1675 660 -1655
rect 360 -1694 362 -1690
rect 398 -1694 400 -1690
rect 324 -1724 326 -1716
rect 620 -1699 622 -1695
rect 658 -1699 660 -1695
rect 584 -1712 586 -1700
rect 491 -1724 493 -1720
rect 529 -1724 531 -1720
rect 324 -1759 326 -1744
rect 360 -1754 362 -1734
rect 398 -1754 400 -1734
rect 455 -1754 457 -1746
rect 360 -1778 362 -1774
rect 398 -1778 400 -1774
rect 324 -1783 326 -1779
rect 455 -1789 457 -1774
rect 491 -1784 493 -1764
rect 529 -1784 531 -1764
rect 749 -1804 751 -1800
rect 787 -1804 789 -1800
rect 491 -1808 493 -1804
rect 529 -1808 531 -1804
rect 455 -1813 457 -1809
rect 713 -1834 715 -1830
rect 360 -1838 362 -1834
rect 398 -1838 400 -1834
rect 324 -1868 326 -1860
rect 713 -1869 715 -1854
rect 749 -1864 751 -1844
rect 787 -1864 789 -1844
rect 324 -1903 326 -1888
rect 360 -1898 362 -1878
rect 398 -1898 400 -1878
rect 749 -1888 751 -1884
rect 787 -1888 789 -1884
rect 713 -1901 715 -1889
rect 360 -1922 362 -1918
rect 398 -1922 400 -1918
rect 324 -1927 326 -1923
rect 360 -1965 362 -1961
rect 398 -1965 400 -1961
rect 324 -1995 326 -1987
rect 491 -1995 493 -1991
rect 529 -1995 531 -1991
rect 324 -2030 326 -2015
rect 360 -2025 362 -2005
rect 398 -2025 400 -2005
rect 455 -2025 457 -2017
rect 626 -2025 628 -2021
rect 664 -2025 666 -2021
rect 360 -2049 362 -2045
rect 398 -2049 400 -2045
rect 324 -2054 326 -2050
rect 455 -2060 457 -2045
rect 491 -2055 493 -2035
rect 529 -2055 531 -2035
rect 590 -2055 592 -2047
rect 491 -2079 493 -2075
rect 529 -2079 531 -2075
rect 455 -2084 457 -2080
rect 590 -2090 592 -2075
rect 626 -2085 628 -2065
rect 664 -2085 666 -2065
rect 360 -2109 362 -2105
rect 398 -2109 400 -2105
rect 324 -2139 326 -2131
rect 626 -2109 628 -2105
rect 664 -2109 666 -2105
rect 590 -2114 592 -2110
rect 324 -2174 326 -2159
rect 360 -2169 362 -2149
rect 398 -2169 400 -2149
rect 360 -2193 362 -2189
rect 398 -2193 400 -2189
rect 324 -2198 326 -2194
<< polycontact >>
rect 373 280 378 285
rect 320 262 325 267
rect 345 239 350 244
rect 405 216 410 221
rect 320 211 325 216
rect 74 118 79 123
rect 143 91 148 96
rect 181 91 186 96
rect 414 99 419 104
rect 452 99 457 104
rect 609 99 614 104
rect 556 81 561 86
rect 378 59 383 64
rect 581 58 586 63
rect 49 46 54 51
rect 111 35 116 40
rect 641 35 646 40
rect 556 30 561 35
rect 58 17 63 22
rect 83 -6 88 -1
rect 272 1 277 6
rect 143 -29 148 -24
rect 58 -34 63 -29
rect 308 -29 313 -24
rect 346 -29 351 -24
rect 74 -172 79 -167
rect 143 -199 148 -194
rect 181 -199 186 -194
rect 491 -191 496 -186
rect 529 -191 534 -186
rect 455 -231 460 -226
rect 49 -244 54 -239
rect 111 -255 116 -250
rect 58 -273 63 -268
rect 83 -296 88 -291
rect 352 -289 357 -284
rect 143 -319 148 -314
rect 58 -324 63 -319
rect 388 -319 393 -314
rect 426 -319 431 -314
rect 611 -313 616 -308
rect 649 -313 654 -308
rect 811 -313 816 -308
rect 758 -331 763 -326
rect 575 -353 580 -348
rect 783 -354 788 -349
rect 843 -377 848 -372
rect 758 -382 763 -377
rect 280 -415 285 -410
rect 316 -445 321 -440
rect 354 -445 359 -440
rect 409 -445 414 -440
rect 445 -475 450 -470
rect 483 -475 488 -470
rect 74 -589 79 -584
rect 143 -616 148 -611
rect 181 -616 186 -611
rect 648 -608 653 -603
rect 686 -608 691 -603
rect 612 -648 617 -643
rect 49 -661 54 -656
rect 111 -672 116 -667
rect 58 -690 63 -685
rect 83 -713 88 -708
rect 304 -706 309 -701
rect 143 -736 148 -731
rect 58 -741 63 -736
rect 340 -736 345 -731
rect 378 -736 383 -731
rect 815 -745 820 -740
rect 853 -745 858 -740
rect 1010 -745 1015 -740
rect 957 -763 962 -758
rect 779 -785 784 -780
rect 982 -786 987 -781
rect 1042 -809 1047 -804
rect 957 -814 962 -809
rect 304 -850 309 -845
rect 340 -880 345 -875
rect 378 -880 383 -875
rect 433 -880 438 -875
rect 469 -910 474 -905
rect 507 -910 512 -905
rect 644 -964 649 -959
rect 682 -964 687 -959
rect 307 -1020 312 -1015
rect 608 -1004 613 -999
rect 343 -1050 348 -1045
rect 381 -1050 386 -1045
rect 438 -1050 443 -1045
rect 474 -1080 479 -1075
rect 512 -1080 517 -1075
rect 307 -1164 312 -1159
rect 343 -1194 348 -1189
rect 381 -1194 386 -1189
rect 74 -1290 79 -1285
rect 143 -1317 148 -1312
rect 181 -1317 186 -1312
rect 49 -1362 54 -1357
rect 111 -1373 116 -1368
rect 58 -1391 63 -1386
rect 83 -1414 88 -1409
rect 316 -1407 321 -1402
rect 143 -1437 148 -1432
rect 58 -1442 63 -1437
rect 506 -1397 511 -1392
rect 544 -1397 549 -1392
rect 352 -1437 357 -1432
rect 390 -1437 395 -1432
rect 470 -1437 475 -1432
rect 855 -1493 860 -1488
rect 893 -1493 898 -1488
rect 316 -1551 321 -1546
rect 819 -1533 824 -1528
rect 352 -1581 357 -1576
rect 390 -1581 395 -1576
rect 445 -1581 450 -1576
rect 481 -1611 486 -1606
rect 519 -1611 524 -1606
rect 615 -1672 620 -1667
rect 653 -1672 658 -1667
rect 319 -1721 324 -1716
rect 579 -1712 584 -1707
rect 355 -1751 360 -1746
rect 393 -1751 398 -1746
rect 450 -1751 455 -1746
rect 486 -1781 491 -1776
rect 524 -1781 529 -1776
rect 319 -1865 324 -1860
rect 744 -1861 749 -1856
rect 782 -1861 787 -1856
rect 355 -1895 360 -1890
rect 393 -1895 398 -1890
rect 708 -1901 713 -1896
rect 319 -1992 324 -1987
rect 355 -2022 360 -2017
rect 393 -2022 398 -2017
rect 450 -2022 455 -2017
rect 486 -2052 491 -2047
rect 524 -2052 529 -2047
rect 585 -2052 590 -2047
rect 621 -2082 626 -2077
rect 659 -2082 664 -2077
rect 319 -2136 324 -2131
rect 355 -2166 360 -2161
rect 393 -2166 398 -2161
<< metal1 >>
rect 395 285 427 288
rect 225 280 373 285
rect 395 281 398 285
rect 402 281 420 285
rect 424 281 427 285
rect 253 274 262 277
rect 253 270 256 274
rect 260 270 262 274
rect 253 267 262 270
rect 320 267 325 280
rect 395 279 427 281
rect 355 275 363 277
rect 355 271 357 275
rect 361 271 363 275
rect 405 273 409 279
rect 355 267 363 271
rect 253 263 268 267
rect 253 252 262 263
rect 348 263 363 267
rect 308 255 328 259
rect 253 248 256 252
rect 260 248 262 252
rect 253 245 262 248
rect 320 244 325 255
rect 355 251 363 263
rect 355 247 357 251
rect 361 247 363 251
rect 373 250 377 252
rect 355 245 363 247
rect 366 246 377 250
rect 381 248 385 252
rect 320 239 345 244
rect 366 235 370 246
rect 381 243 394 248
rect 381 240 385 243
rect 234 230 370 235
rect 253 223 262 226
rect 253 219 256 223
rect 260 219 262 223
rect 253 216 262 219
rect 320 216 325 230
rect 355 224 363 226
rect 355 220 357 224
rect 361 220 363 224
rect 355 216 363 220
rect 253 212 268 216
rect 253 201 262 212
rect 348 212 363 216
rect 308 204 328 208
rect 253 197 256 201
rect 260 197 262 201
rect 253 194 262 197
rect 320 189 325 204
rect 355 200 363 212
rect 355 196 357 200
rect 361 196 363 200
rect 355 194 363 196
rect 389 221 394 243
rect 413 221 417 233
rect 373 189 377 220
rect 389 216 405 221
rect 413 216 427 221
rect 413 213 417 216
rect 320 184 377 189
rect 405 186 409 193
rect 395 184 427 186
rect 395 180 397 184
rect 401 180 421 184
rect 425 180 427 184
rect 395 178 427 180
rect 378 168 474 171
rect 378 164 407 168
rect 411 164 467 168
rect 471 164 474 168
rect 133 160 165 163
rect 133 156 136 160
rect 140 156 158 160
rect 162 156 165 160
rect 133 154 165 156
rect 171 160 203 163
rect 171 156 174 160
rect 178 156 196 160
rect 200 156 203 160
rect 171 154 203 156
rect 378 162 474 164
rect 143 148 147 154
rect 181 148 185 154
rect -22 95 58 100
rect -22 -10 -17 95
rect -9 29 0 32
rect -9 25 -6 29
rect -2 25 0 29
rect -9 22 0 25
rect -9 18 6 22
rect -9 7 0 18
rect 49 14 54 46
rect 74 40 79 118
rect 111 100 115 101
rect 95 95 115 100
rect 119 96 123 101
rect 151 96 155 108
rect 189 96 193 108
rect 378 126 382 162
rect 414 156 418 162
rect 452 156 456 162
rect 386 104 390 106
rect 422 104 426 116
rect 460 104 464 116
rect 631 104 663 107
rect 386 99 414 104
rect 422 99 452 104
rect 460 99 609 104
rect 631 100 634 104
rect 638 100 656 104
rect 660 100 663 104
rect 119 91 143 96
rect 151 91 181 96
rect 189 91 238 96
rect 243 91 383 96
rect 386 91 390 99
rect 422 96 426 99
rect 460 96 464 99
rect 119 89 123 91
rect 151 88 155 91
rect 189 88 193 91
rect 111 67 115 69
rect 102 66 115 67
rect 102 62 103 66
rect 107 62 115 66
rect 102 61 115 62
rect 489 93 498 96
rect 489 89 492 93
rect 496 89 498 93
rect 489 86 498 89
rect 556 86 561 99
rect 631 98 663 100
rect 591 94 599 96
rect 591 90 593 94
rect 597 90 599 94
rect 641 92 645 98
rect 591 86 599 90
rect 489 82 504 86
rect 143 61 147 68
rect 181 61 185 68
rect 133 59 165 61
rect 133 55 135 59
rect 139 55 159 59
rect 163 55 165 59
rect 133 53 165 55
rect 171 59 203 61
rect 171 55 173 59
rect 177 55 197 59
rect 201 55 203 59
rect 171 53 203 55
rect 414 62 418 76
rect 452 62 456 76
rect 489 71 498 82
rect 584 82 599 86
rect 544 74 564 78
rect 489 67 492 71
rect 496 67 498 71
rect 489 64 498 67
rect 556 63 561 74
rect 591 70 599 82
rect 591 66 593 70
rect 597 66 599 70
rect 609 69 613 71
rect 591 64 599 66
rect 602 65 613 69
rect 617 67 621 71
rect 133 40 165 43
rect 58 35 111 40
rect 133 36 136 40
rect 140 36 158 40
rect 162 36 165 40
rect 58 22 63 35
rect 133 34 165 36
rect 298 40 368 43
rect 298 36 301 40
rect 305 36 361 40
rect 365 36 368 40
rect 298 34 368 36
rect 93 30 101 32
rect 93 26 95 30
rect 99 26 101 30
rect 143 28 147 34
rect 308 28 312 34
rect 346 28 350 34
rect 93 22 101 26
rect 86 18 101 22
rect 46 10 66 14
rect -9 3 -6 7
rect -2 3 0 7
rect -9 0 0 3
rect 58 -1 63 10
rect 93 6 101 18
rect 93 2 95 6
rect 99 2 101 6
rect 111 5 115 7
rect 93 0 101 2
rect 104 1 115 5
rect 119 3 123 7
rect 58 -6 83 -1
rect 104 -10 108 1
rect 119 -2 132 3
rect 119 -5 123 -2
rect -22 -15 108 -10
rect -9 -22 0 -19
rect -9 -26 -6 -22
rect -2 -26 0 -22
rect -9 -29 0 -26
rect 58 -29 63 -15
rect 93 -21 101 -19
rect 93 -25 95 -21
rect 99 -25 101 -21
rect 93 -29 101 -25
rect -9 -33 6 -29
rect -9 -44 0 -33
rect 86 -33 101 -29
rect 46 -41 66 -37
rect -9 -48 -6 -44
rect -2 -48 0 -44
rect -9 -51 0 -48
rect 58 -56 63 -41
rect 93 -45 101 -33
rect 93 -49 95 -45
rect 99 -49 101 -45
rect 93 -51 101 -49
rect 127 -24 132 -2
rect 234 1 272 6
rect 151 -24 155 -12
rect 272 -24 276 -22
rect 111 -56 115 -25
rect 127 -29 143 -24
rect 151 -29 220 -24
rect 225 -29 276 -24
rect 280 -24 284 -22
rect 316 -24 320 -12
rect 354 -24 358 -12
rect 378 -24 383 59
rect 404 60 474 62
rect 404 56 406 60
rect 410 56 468 60
rect 472 56 474 60
rect 556 58 581 63
rect 404 54 474 56
rect 602 54 606 65
rect 617 62 630 67
rect 617 59 621 62
rect 494 49 606 54
rect 489 42 498 45
rect 489 38 492 42
rect 496 38 498 42
rect 489 35 498 38
rect 556 35 561 49
rect 591 43 599 45
rect 591 39 593 43
rect 597 39 599 43
rect 591 35 599 39
rect 489 31 504 35
rect 489 20 498 31
rect 584 31 599 35
rect 544 23 564 27
rect 489 16 492 20
rect 496 16 498 20
rect 489 13 498 16
rect 556 8 561 23
rect 591 19 599 31
rect 591 15 593 19
rect 597 15 599 19
rect 591 13 599 15
rect 625 40 630 62
rect 649 40 653 52
rect 609 8 613 39
rect 625 35 641 40
rect 649 35 663 40
rect 649 32 653 35
rect 556 3 613 8
rect 641 5 645 12
rect 631 3 663 5
rect 631 -1 633 3
rect 637 -1 657 3
rect 661 -1 663 3
rect 631 -3 663 -1
rect 280 -29 308 -24
rect 316 -29 346 -24
rect 354 -29 383 -24
rect 151 -32 155 -29
rect 58 -61 115 -56
rect 280 -37 284 -29
rect 316 -32 320 -29
rect 354 -32 358 -29
rect 143 -59 147 -52
rect 133 -61 165 -59
rect 133 -65 135 -61
rect 139 -65 159 -61
rect 163 -65 165 -61
rect 133 -67 165 -65
rect 272 -66 276 -57
rect 308 -66 312 -52
rect 346 -66 350 -52
rect 262 -68 368 -66
rect 262 -72 264 -68
rect 268 -72 362 -68
rect 366 -72 368 -68
rect 262 -74 368 -72
rect 252 -86 464 -81
rect 455 -122 551 -119
rect 455 -126 484 -122
rect 488 -126 544 -122
rect 548 -126 551 -122
rect 133 -130 165 -127
rect 133 -134 136 -130
rect 140 -134 158 -130
rect 162 -134 165 -130
rect 133 -136 165 -134
rect 171 -130 203 -127
rect 171 -134 174 -130
rect 178 -134 196 -130
rect 200 -134 203 -130
rect 171 -136 203 -134
rect 455 -128 551 -126
rect 143 -142 147 -136
rect 181 -142 185 -136
rect -22 -195 58 -190
rect -22 -300 -17 -195
rect -9 -261 0 -258
rect -9 -265 -6 -261
rect -2 -265 0 -261
rect -9 -268 0 -265
rect -9 -272 6 -268
rect -9 -283 0 -272
rect 49 -276 54 -244
rect 74 -250 79 -172
rect 111 -190 115 -189
rect 95 -195 115 -190
rect 119 -194 123 -189
rect 151 -194 155 -182
rect 189 -194 193 -182
rect 455 -164 459 -128
rect 491 -134 495 -128
rect 529 -134 533 -128
rect 463 -186 467 -184
rect 499 -186 503 -174
rect 537 -186 541 -174
rect 463 -191 491 -186
rect 499 -191 529 -186
rect 537 -191 560 -186
rect 119 -199 143 -194
rect 151 -199 181 -194
rect 189 -199 256 -194
rect 261 -199 460 -194
rect 463 -199 467 -191
rect 499 -194 503 -191
rect 537 -194 541 -191
rect 119 -201 123 -199
rect 151 -202 155 -199
rect 189 -202 193 -199
rect 111 -223 115 -221
rect 102 -224 115 -223
rect 102 -228 103 -224
rect 107 -228 115 -224
rect 102 -229 115 -228
rect 143 -229 147 -222
rect 181 -229 185 -222
rect 133 -231 165 -229
rect 133 -235 135 -231
rect 139 -235 159 -231
rect 163 -235 165 -231
rect 133 -237 165 -235
rect 171 -231 203 -229
rect 171 -235 173 -231
rect 177 -235 197 -231
rect 201 -235 203 -231
rect 171 -237 203 -235
rect 491 -228 495 -214
rect 529 -228 533 -214
rect 133 -250 165 -247
rect 58 -255 111 -250
rect 133 -254 136 -250
rect 140 -254 158 -250
rect 162 -254 165 -250
rect 58 -268 63 -255
rect 133 -256 165 -254
rect 378 -250 448 -247
rect 378 -254 381 -250
rect 385 -254 441 -250
rect 445 -254 448 -250
rect 378 -256 448 -254
rect 93 -260 101 -258
rect 93 -264 95 -260
rect 99 -264 101 -260
rect 143 -262 147 -256
rect 388 -262 392 -256
rect 426 -262 430 -256
rect 93 -268 101 -264
rect 86 -272 101 -268
rect 46 -280 66 -276
rect -9 -287 -6 -283
rect -2 -287 0 -283
rect -9 -290 0 -287
rect 58 -291 63 -280
rect 93 -284 101 -272
rect 93 -288 95 -284
rect 99 -288 101 -284
rect 111 -285 115 -283
rect 93 -290 101 -288
rect 104 -289 115 -285
rect 119 -287 123 -283
rect 58 -296 83 -291
rect 104 -300 108 -289
rect 119 -292 132 -287
rect 119 -295 123 -292
rect -22 -305 108 -300
rect -9 -312 0 -309
rect -9 -316 -6 -312
rect -2 -316 0 -312
rect -9 -319 0 -316
rect 58 -319 63 -305
rect 93 -311 101 -309
rect 93 -315 95 -311
rect 99 -315 101 -311
rect 93 -319 101 -315
rect -9 -323 6 -319
rect -9 -334 0 -323
rect 86 -323 101 -319
rect 46 -331 66 -327
rect -9 -338 -6 -334
rect -2 -338 0 -334
rect -9 -341 0 -338
rect 58 -346 63 -331
rect 93 -335 101 -323
rect 93 -339 95 -335
rect 99 -339 101 -335
rect 93 -341 101 -339
rect 127 -314 132 -292
rect 243 -289 352 -284
rect 151 -314 155 -302
rect 352 -314 356 -312
rect 111 -346 115 -315
rect 127 -319 143 -314
rect 151 -319 247 -314
rect 252 -319 356 -314
rect 360 -314 364 -312
rect 396 -314 400 -302
rect 434 -314 438 -302
rect 455 -314 460 -231
rect 481 -230 551 -228
rect 481 -234 483 -230
rect 487 -234 545 -230
rect 549 -234 551 -230
rect 481 -236 551 -234
rect 360 -319 388 -314
rect 396 -319 426 -314
rect 434 -319 460 -314
rect 555 -316 560 -191
rect 575 -244 671 -241
rect 575 -248 604 -244
rect 608 -248 664 -244
rect 668 -248 671 -244
rect 575 -250 671 -248
rect 575 -286 579 -250
rect 611 -256 615 -250
rect 649 -256 653 -250
rect 583 -308 587 -306
rect 619 -308 623 -296
rect 657 -308 661 -296
rect 833 -308 865 -305
rect 583 -313 611 -308
rect 619 -313 649 -308
rect 657 -313 811 -308
rect 833 -312 836 -308
rect 840 -312 858 -308
rect 862 -312 865 -308
rect 151 -322 155 -319
rect 58 -351 115 -346
rect 360 -327 364 -319
rect 396 -322 400 -319
rect 434 -322 438 -319
rect 555 -321 580 -316
rect 583 -321 587 -313
rect 619 -316 623 -313
rect 657 -316 661 -313
rect 143 -349 147 -342
rect 691 -319 700 -316
rect 691 -323 694 -319
rect 698 -323 700 -319
rect 691 -326 700 -323
rect 758 -326 763 -313
rect 833 -314 865 -312
rect 793 -318 801 -316
rect 793 -322 795 -318
rect 799 -322 801 -318
rect 843 -320 847 -314
rect 793 -326 801 -322
rect 691 -330 706 -326
rect 133 -351 165 -349
rect 133 -355 135 -351
rect 139 -355 159 -351
rect 163 -355 165 -351
rect 133 -357 165 -355
rect 352 -356 356 -347
rect 388 -356 392 -342
rect 426 -356 430 -342
rect 565 -353 575 -348
rect 611 -350 615 -336
rect 649 -350 653 -336
rect 691 -341 700 -330
rect 786 -330 801 -326
rect 746 -338 766 -334
rect 691 -345 694 -341
rect 698 -345 700 -341
rect 691 -348 700 -345
rect 758 -349 763 -338
rect 793 -342 801 -330
rect 793 -346 795 -342
rect 799 -346 801 -342
rect 811 -343 815 -341
rect 793 -348 801 -346
rect 804 -347 815 -343
rect 819 -345 823 -341
rect 601 -352 671 -350
rect 342 -358 448 -356
rect 342 -362 344 -358
rect 348 -362 442 -358
rect 446 -362 448 -358
rect 342 -364 448 -362
rect 306 -376 376 -373
rect 306 -380 309 -376
rect 313 -380 369 -376
rect 373 -380 376 -376
rect 306 -382 376 -380
rect 316 -388 320 -382
rect 354 -388 358 -382
rect 225 -415 280 -410
rect 280 -440 284 -438
rect 234 -445 284 -440
rect 435 -406 505 -403
rect 435 -410 438 -406
rect 442 -410 498 -406
rect 502 -410 505 -406
rect 435 -412 505 -410
rect 288 -440 292 -438
rect 324 -440 328 -428
rect 362 -440 366 -428
rect 445 -418 449 -412
rect 483 -418 487 -412
rect 288 -445 316 -440
rect 324 -445 354 -440
rect 362 -445 409 -440
rect 288 -453 292 -445
rect 324 -448 328 -445
rect 362 -448 366 -445
rect 280 -482 284 -473
rect 316 -482 320 -468
rect 354 -482 358 -468
rect 409 -470 413 -468
rect 389 -475 413 -470
rect 417 -470 421 -468
rect 453 -470 457 -458
rect 491 -470 495 -458
rect 565 -470 570 -353
rect 601 -356 603 -352
rect 607 -356 665 -352
rect 669 -356 671 -352
rect 758 -354 783 -349
rect 601 -358 671 -356
rect 804 -358 808 -347
rect 819 -350 832 -345
rect 819 -353 823 -350
rect 696 -363 808 -358
rect 691 -370 700 -367
rect 691 -374 694 -370
rect 698 -374 700 -370
rect 691 -377 700 -374
rect 758 -377 763 -363
rect 793 -369 801 -367
rect 793 -373 795 -369
rect 799 -373 801 -369
rect 793 -377 801 -373
rect 691 -381 706 -377
rect 691 -392 700 -381
rect 786 -381 801 -377
rect 746 -389 766 -385
rect 691 -396 694 -392
rect 698 -396 700 -392
rect 691 -399 700 -396
rect 758 -404 763 -389
rect 793 -393 801 -381
rect 793 -397 795 -393
rect 799 -397 801 -393
rect 793 -399 801 -397
rect 827 -372 832 -350
rect 851 -372 855 -360
rect 811 -404 815 -373
rect 827 -377 843 -372
rect 851 -377 865 -372
rect 851 -380 855 -377
rect 758 -409 815 -404
rect 843 -407 847 -400
rect 833 -409 865 -407
rect 833 -413 835 -409
rect 839 -413 859 -409
rect 863 -413 865 -409
rect 833 -415 865 -413
rect 417 -475 445 -470
rect 453 -475 483 -470
rect 491 -475 570 -470
rect 270 -484 376 -482
rect 270 -488 272 -484
rect 276 -488 370 -484
rect 374 -488 376 -484
rect 270 -490 376 -488
rect 389 -505 395 -475
rect 417 -483 421 -475
rect 453 -478 457 -475
rect 491 -478 495 -475
rect 252 -511 395 -505
rect 409 -512 413 -503
rect 445 -512 449 -498
rect 483 -512 487 -498
rect 399 -514 505 -512
rect 399 -518 401 -514
rect 405 -518 499 -514
rect 503 -518 505 -514
rect 399 -520 505 -518
rect 270 -533 645 -528
rect 612 -539 708 -536
rect 612 -543 641 -539
rect 645 -543 701 -539
rect 705 -543 708 -539
rect 133 -547 165 -544
rect 133 -551 136 -547
rect 140 -551 158 -547
rect 162 -551 165 -547
rect 133 -553 165 -551
rect 171 -547 203 -544
rect 171 -551 174 -547
rect 178 -551 196 -547
rect 200 -551 203 -547
rect 171 -553 203 -551
rect 612 -545 708 -543
rect 143 -559 147 -553
rect 181 -559 185 -553
rect -22 -612 58 -607
rect -22 -717 -17 -612
rect -9 -678 0 -675
rect -9 -682 -6 -678
rect -2 -682 0 -678
rect -9 -685 0 -682
rect -9 -689 6 -685
rect -9 -700 0 -689
rect 49 -693 54 -661
rect 74 -667 79 -589
rect 111 -607 115 -606
rect 95 -612 115 -607
rect 119 -611 123 -606
rect 151 -611 155 -599
rect 189 -611 193 -599
rect 612 -581 616 -545
rect 648 -551 652 -545
rect 686 -551 690 -545
rect 620 -603 624 -601
rect 656 -603 660 -591
rect 694 -603 698 -591
rect 620 -608 648 -603
rect 656 -608 686 -603
rect 694 -608 766 -603
rect 119 -616 143 -611
rect 151 -616 181 -611
rect 189 -616 274 -611
rect 279 -616 617 -611
rect 620 -616 624 -608
rect 656 -611 660 -608
rect 694 -611 698 -608
rect 119 -618 123 -616
rect 151 -619 155 -616
rect 189 -619 193 -616
rect 111 -640 115 -638
rect 102 -641 115 -640
rect 102 -645 103 -641
rect 107 -645 115 -641
rect 102 -646 115 -645
rect 143 -646 147 -639
rect 181 -646 185 -639
rect 133 -648 165 -646
rect 133 -652 135 -648
rect 139 -652 159 -648
rect 163 -652 165 -648
rect 133 -654 165 -652
rect 171 -648 203 -646
rect 171 -652 173 -648
rect 177 -652 197 -648
rect 201 -652 203 -648
rect 171 -654 203 -652
rect 602 -648 612 -643
rect 648 -645 652 -631
rect 686 -645 690 -631
rect 638 -647 708 -645
rect 133 -667 165 -664
rect 58 -672 111 -667
rect 133 -671 136 -667
rect 140 -671 158 -667
rect 162 -671 165 -667
rect 58 -685 63 -672
rect 133 -673 165 -671
rect 330 -667 400 -664
rect 330 -671 333 -667
rect 337 -671 393 -667
rect 397 -671 400 -667
rect 330 -673 400 -671
rect 93 -677 101 -675
rect 93 -681 95 -677
rect 99 -681 101 -677
rect 143 -679 147 -673
rect 340 -679 344 -673
rect 378 -679 382 -673
rect 93 -685 101 -681
rect 86 -689 101 -685
rect 46 -697 66 -693
rect -9 -704 -6 -700
rect -2 -704 0 -700
rect -9 -707 0 -704
rect 58 -708 63 -697
rect 93 -701 101 -689
rect 93 -705 95 -701
rect 99 -705 101 -701
rect 111 -702 115 -700
rect 93 -707 101 -705
rect 104 -706 115 -702
rect 119 -704 123 -700
rect 58 -713 83 -708
rect 104 -717 108 -706
rect 119 -709 132 -704
rect 119 -712 123 -709
rect -22 -722 108 -717
rect -9 -729 0 -726
rect -9 -733 -6 -729
rect -2 -733 0 -729
rect -9 -736 0 -733
rect 58 -736 63 -722
rect 93 -728 101 -726
rect 93 -732 95 -728
rect 99 -732 101 -728
rect 93 -736 101 -732
rect -9 -740 6 -736
rect -9 -751 0 -740
rect 86 -740 101 -736
rect 46 -748 66 -744
rect -9 -755 -6 -751
rect -2 -755 0 -751
rect -9 -758 0 -755
rect 58 -763 63 -748
rect 93 -752 101 -740
rect 93 -756 95 -752
rect 99 -756 101 -752
rect 93 -758 101 -756
rect 127 -731 132 -709
rect 261 -706 304 -701
rect 151 -731 155 -719
rect 304 -731 308 -729
rect 111 -763 115 -732
rect 127 -736 143 -731
rect 151 -736 265 -731
rect 270 -736 308 -731
rect 312 -731 316 -729
rect 348 -731 352 -719
rect 386 -731 390 -719
rect 602 -731 607 -648
rect 638 -651 640 -647
rect 644 -651 702 -647
rect 706 -651 708 -647
rect 638 -653 708 -651
rect 312 -736 340 -731
rect 348 -736 378 -731
rect 386 -736 607 -731
rect 151 -739 155 -736
rect 58 -768 115 -763
rect 312 -744 316 -736
rect 348 -739 352 -736
rect 386 -739 390 -736
rect 143 -766 147 -759
rect 761 -748 766 -608
rect 779 -676 875 -673
rect 779 -680 808 -676
rect 812 -680 868 -676
rect 872 -680 875 -676
rect 779 -682 875 -680
rect 779 -718 783 -682
rect 815 -688 819 -682
rect 853 -688 857 -682
rect 787 -740 791 -738
rect 823 -740 827 -728
rect 861 -740 865 -728
rect 1032 -740 1064 -737
rect 787 -745 815 -740
rect 823 -745 853 -740
rect 861 -745 1010 -740
rect 1032 -744 1035 -740
rect 1039 -744 1057 -740
rect 1061 -744 1064 -740
rect 761 -753 784 -748
rect 787 -753 791 -745
rect 823 -748 827 -745
rect 861 -748 865 -745
rect 133 -768 165 -766
rect 133 -772 135 -768
rect 139 -772 159 -768
rect 163 -772 165 -768
rect 133 -774 165 -772
rect 304 -773 308 -764
rect 340 -773 344 -759
rect 378 -773 382 -759
rect 890 -751 899 -748
rect 890 -755 893 -751
rect 897 -755 899 -751
rect 890 -758 899 -755
rect 957 -758 962 -745
rect 1032 -746 1064 -744
rect 992 -750 1000 -748
rect 992 -754 994 -750
rect 998 -754 1000 -750
rect 1042 -752 1046 -746
rect 992 -758 1000 -754
rect 890 -762 905 -758
rect 294 -775 400 -773
rect 294 -779 296 -775
rect 300 -779 394 -775
rect 398 -779 400 -775
rect 294 -781 400 -779
rect 761 -785 779 -780
rect 815 -782 819 -768
rect 853 -782 857 -768
rect 890 -773 899 -762
rect 985 -762 1000 -758
rect 945 -770 965 -766
rect 890 -777 893 -773
rect 897 -777 899 -773
rect 890 -780 899 -777
rect 957 -781 962 -770
rect 992 -774 1000 -762
rect 992 -778 994 -774
rect 998 -778 1000 -774
rect 1010 -775 1014 -773
rect 992 -780 1000 -778
rect 1003 -779 1014 -775
rect 1018 -777 1022 -773
rect 805 -784 875 -782
rect 330 -811 400 -808
rect 330 -815 333 -811
rect 337 -815 393 -811
rect 397 -815 400 -811
rect 330 -817 400 -815
rect 340 -823 344 -817
rect 378 -823 382 -817
rect 243 -850 304 -845
rect 304 -875 308 -873
rect 252 -880 308 -875
rect 459 -841 529 -838
rect 459 -845 462 -841
rect 466 -845 522 -841
rect 526 -845 529 -841
rect 459 -847 529 -845
rect 312 -875 316 -873
rect 348 -875 352 -863
rect 386 -875 390 -863
rect 469 -853 473 -847
rect 507 -853 511 -847
rect 312 -880 340 -875
rect 348 -880 378 -875
rect 386 -880 433 -875
rect 312 -888 316 -880
rect 348 -883 352 -880
rect 386 -883 390 -880
rect 304 -917 308 -908
rect 340 -917 344 -903
rect 378 -917 382 -903
rect 433 -905 437 -903
rect 413 -910 437 -905
rect 441 -905 445 -903
rect 477 -905 481 -893
rect 515 -905 519 -893
rect 608 -895 704 -892
rect 608 -899 637 -895
rect 641 -899 697 -895
rect 701 -899 704 -895
rect 608 -901 704 -899
rect 441 -910 469 -905
rect 477 -910 507 -905
rect 515 -910 581 -905
rect 294 -919 400 -917
rect 294 -923 296 -919
rect 300 -923 394 -919
rect 398 -923 400 -919
rect 294 -925 400 -923
rect 413 -940 419 -910
rect 441 -918 445 -910
rect 477 -913 481 -910
rect 515 -913 519 -910
rect 270 -945 419 -940
rect 433 -947 437 -938
rect 469 -947 473 -933
rect 507 -947 511 -933
rect 423 -949 529 -947
rect 423 -953 425 -949
rect 429 -953 523 -949
rect 527 -953 529 -949
rect 423 -955 529 -953
rect 576 -967 581 -910
rect 608 -937 612 -901
rect 644 -907 648 -901
rect 682 -907 686 -901
rect 616 -959 620 -957
rect 652 -959 656 -947
rect 690 -959 694 -947
rect 761 -959 766 -785
rect 805 -788 807 -784
rect 811 -788 869 -784
rect 873 -788 875 -784
rect 957 -786 982 -781
rect 805 -790 875 -788
rect 1003 -790 1007 -779
rect 1018 -782 1031 -777
rect 1018 -785 1022 -782
rect 895 -795 1007 -790
rect 890 -802 899 -799
rect 890 -806 893 -802
rect 897 -806 899 -802
rect 890 -809 899 -806
rect 957 -809 962 -795
rect 992 -801 1000 -799
rect 992 -805 994 -801
rect 998 -805 1000 -801
rect 992 -809 1000 -805
rect 890 -813 905 -809
rect 890 -824 899 -813
rect 985 -813 1000 -809
rect 945 -821 965 -817
rect 890 -828 893 -824
rect 897 -828 899 -824
rect 890 -831 899 -828
rect 957 -836 962 -821
rect 992 -825 1000 -813
rect 992 -829 994 -825
rect 998 -829 1000 -825
rect 992 -831 1000 -829
rect 1026 -804 1031 -782
rect 1050 -804 1054 -792
rect 1010 -836 1014 -805
rect 1026 -809 1042 -804
rect 1050 -809 1064 -804
rect 1050 -812 1054 -809
rect 957 -841 1014 -836
rect 1042 -839 1046 -832
rect 1032 -841 1064 -839
rect 1032 -845 1034 -841
rect 1038 -845 1058 -841
rect 1062 -845 1064 -841
rect 1032 -847 1064 -845
rect 616 -964 644 -959
rect 652 -964 682 -959
rect 690 -964 766 -959
rect 576 -972 613 -967
rect 616 -972 620 -964
rect 652 -967 656 -964
rect 690 -967 694 -964
rect 333 -981 403 -978
rect 333 -985 336 -981
rect 340 -985 396 -981
rect 400 -985 403 -981
rect 333 -987 403 -985
rect 343 -993 347 -987
rect 381 -993 385 -987
rect 225 -1020 307 -1015
rect 307 -1045 311 -1043
rect 234 -1050 311 -1045
rect 598 -1004 608 -999
rect 644 -1001 648 -987
rect 682 -1001 686 -987
rect 634 -1003 704 -1001
rect 464 -1011 534 -1008
rect 464 -1015 467 -1011
rect 471 -1015 527 -1011
rect 531 -1015 534 -1011
rect 464 -1017 534 -1015
rect 315 -1045 319 -1043
rect 351 -1045 355 -1033
rect 389 -1045 393 -1033
rect 474 -1023 478 -1017
rect 512 -1023 516 -1017
rect 315 -1050 343 -1045
rect 351 -1050 381 -1045
rect 389 -1050 438 -1045
rect 315 -1058 319 -1050
rect 351 -1053 355 -1050
rect 389 -1053 393 -1050
rect 307 -1087 311 -1078
rect 343 -1087 347 -1073
rect 381 -1087 385 -1073
rect 438 -1075 442 -1073
rect 408 -1080 442 -1075
rect 446 -1075 450 -1073
rect 482 -1075 486 -1063
rect 520 -1075 524 -1063
rect 598 -1075 604 -1004
rect 634 -1007 636 -1003
rect 640 -1007 698 -1003
rect 702 -1007 704 -1003
rect 634 -1009 704 -1007
rect 446 -1080 474 -1075
rect 482 -1080 512 -1075
rect 520 -1080 604 -1075
rect 297 -1089 403 -1087
rect 297 -1093 299 -1089
rect 303 -1093 397 -1089
rect 401 -1093 403 -1089
rect 297 -1095 403 -1093
rect 333 -1125 403 -1122
rect 333 -1129 336 -1125
rect 340 -1129 396 -1125
rect 400 -1129 403 -1125
rect 333 -1131 403 -1129
rect 343 -1137 347 -1131
rect 381 -1137 385 -1131
rect 252 -1164 307 -1159
rect 307 -1189 311 -1187
rect 270 -1194 311 -1189
rect 315 -1189 319 -1187
rect 351 -1189 355 -1177
rect 389 -1189 393 -1177
rect 408 -1189 413 -1080
rect 446 -1088 450 -1080
rect 482 -1083 486 -1080
rect 520 -1083 524 -1080
rect 438 -1117 442 -1108
rect 474 -1117 478 -1103
rect 512 -1117 516 -1103
rect 428 -1119 534 -1117
rect 428 -1123 430 -1119
rect 434 -1123 528 -1119
rect 532 -1123 534 -1119
rect 428 -1125 534 -1123
rect 315 -1194 343 -1189
rect 351 -1194 381 -1189
rect 389 -1194 413 -1189
rect 315 -1202 319 -1194
rect 351 -1197 355 -1194
rect 389 -1197 393 -1194
rect 307 -1231 311 -1222
rect 343 -1231 347 -1217
rect 381 -1231 385 -1217
rect 297 -1233 403 -1231
rect 297 -1237 299 -1233
rect 303 -1237 397 -1233
rect 401 -1237 403 -1233
rect 297 -1239 403 -1237
rect 133 -1248 165 -1245
rect 133 -1252 136 -1248
rect 140 -1252 158 -1248
rect 162 -1252 165 -1248
rect 133 -1254 165 -1252
rect 171 -1248 203 -1245
rect 171 -1252 174 -1248
rect 178 -1252 196 -1248
rect 200 -1252 203 -1248
rect 288 -1249 853 -1244
rect 171 -1254 203 -1252
rect 143 -1260 147 -1254
rect 181 -1260 185 -1254
rect -22 -1313 58 -1308
rect -22 -1418 -17 -1313
rect -9 -1379 0 -1376
rect -9 -1383 -6 -1379
rect -2 -1383 0 -1379
rect -9 -1386 0 -1383
rect -9 -1390 6 -1386
rect -9 -1401 0 -1390
rect 49 -1394 54 -1362
rect 74 -1368 79 -1290
rect 111 -1308 115 -1307
rect 95 -1313 115 -1308
rect 119 -1312 123 -1307
rect 151 -1312 155 -1300
rect 189 -1312 193 -1300
rect 119 -1317 143 -1312
rect 151 -1317 181 -1312
rect 189 -1317 465 -1312
rect 119 -1319 123 -1317
rect 151 -1320 155 -1317
rect 189 -1320 193 -1317
rect 111 -1341 115 -1339
rect 102 -1342 115 -1341
rect 102 -1346 103 -1342
rect 107 -1346 115 -1342
rect 102 -1347 115 -1346
rect 143 -1347 147 -1340
rect 181 -1347 185 -1340
rect 133 -1349 165 -1347
rect 133 -1353 135 -1349
rect 139 -1353 159 -1349
rect 163 -1353 165 -1349
rect 133 -1355 165 -1353
rect 171 -1349 203 -1347
rect 171 -1353 173 -1349
rect 177 -1353 197 -1349
rect 201 -1353 203 -1349
rect 171 -1355 203 -1353
rect 133 -1368 165 -1365
rect 58 -1373 111 -1368
rect 133 -1372 136 -1368
rect 140 -1372 158 -1368
rect 162 -1372 165 -1368
rect 58 -1386 63 -1373
rect 133 -1374 165 -1372
rect 342 -1368 412 -1365
rect 342 -1372 345 -1368
rect 349 -1372 405 -1368
rect 409 -1372 412 -1368
rect 342 -1374 412 -1372
rect 93 -1378 101 -1376
rect 93 -1382 95 -1378
rect 99 -1382 101 -1378
rect 143 -1380 147 -1374
rect 352 -1380 356 -1374
rect 390 -1380 394 -1374
rect 93 -1386 101 -1382
rect 86 -1390 101 -1386
rect 46 -1398 66 -1394
rect -9 -1405 -6 -1401
rect -2 -1405 0 -1401
rect -9 -1408 0 -1405
rect 58 -1409 63 -1398
rect 93 -1402 101 -1390
rect 93 -1406 95 -1402
rect 99 -1406 101 -1402
rect 111 -1403 115 -1401
rect 93 -1408 101 -1406
rect 104 -1407 115 -1403
rect 119 -1405 123 -1401
rect 58 -1414 83 -1409
rect 104 -1418 108 -1407
rect 119 -1410 132 -1405
rect 119 -1413 123 -1410
rect -22 -1423 108 -1418
rect -9 -1430 0 -1427
rect -9 -1434 -6 -1430
rect -2 -1434 0 -1430
rect -9 -1437 0 -1434
rect 58 -1437 63 -1423
rect 93 -1429 101 -1427
rect 93 -1433 95 -1429
rect 99 -1433 101 -1429
rect 93 -1437 101 -1433
rect -9 -1441 6 -1437
rect -9 -1452 0 -1441
rect 86 -1441 101 -1437
rect 46 -1449 66 -1445
rect -9 -1456 -6 -1452
rect -2 -1456 0 -1452
rect -9 -1459 0 -1456
rect 58 -1464 63 -1449
rect 93 -1453 101 -1441
rect 93 -1457 95 -1453
rect 99 -1457 101 -1453
rect 93 -1459 101 -1457
rect 127 -1432 132 -1410
rect 279 -1407 316 -1402
rect 151 -1432 155 -1420
rect 316 -1432 320 -1430
rect 111 -1464 115 -1433
rect 127 -1437 143 -1432
rect 151 -1437 283 -1432
rect 288 -1437 320 -1432
rect 460 -1400 465 -1317
rect 470 -1328 566 -1325
rect 470 -1332 499 -1328
rect 503 -1332 559 -1328
rect 563 -1332 566 -1328
rect 470 -1334 566 -1332
rect 470 -1370 474 -1334
rect 506 -1340 510 -1334
rect 544 -1340 548 -1334
rect 478 -1392 482 -1390
rect 514 -1392 518 -1380
rect 552 -1392 556 -1380
rect 478 -1397 506 -1392
rect 514 -1397 544 -1392
rect 552 -1397 809 -1392
rect 460 -1405 475 -1400
rect 478 -1405 482 -1397
rect 514 -1400 518 -1397
rect 552 -1400 556 -1397
rect 324 -1432 328 -1430
rect 360 -1432 364 -1420
rect 398 -1432 402 -1420
rect 324 -1437 352 -1432
rect 360 -1437 390 -1432
rect 398 -1437 470 -1432
rect 506 -1434 510 -1420
rect 544 -1434 548 -1420
rect 496 -1436 566 -1434
rect 151 -1440 155 -1437
rect 58 -1469 115 -1464
rect 324 -1445 328 -1437
rect 360 -1440 364 -1437
rect 398 -1440 402 -1437
rect 143 -1467 147 -1460
rect 496 -1440 498 -1436
rect 502 -1440 560 -1436
rect 564 -1440 566 -1436
rect 496 -1442 566 -1440
rect 133 -1469 165 -1467
rect 133 -1473 135 -1469
rect 139 -1473 159 -1469
rect 163 -1473 165 -1469
rect 133 -1475 165 -1473
rect 316 -1474 320 -1465
rect 352 -1474 356 -1460
rect 390 -1474 394 -1460
rect 306 -1476 412 -1474
rect 306 -1480 308 -1476
rect 312 -1480 406 -1476
rect 410 -1480 412 -1476
rect 306 -1482 412 -1480
rect 804 -1496 809 -1397
rect 819 -1424 915 -1421
rect 819 -1428 848 -1424
rect 852 -1428 908 -1424
rect 912 -1428 915 -1424
rect 819 -1430 915 -1428
rect 819 -1466 823 -1430
rect 855 -1436 859 -1430
rect 893 -1436 897 -1430
rect 827 -1488 831 -1486
rect 863 -1488 867 -1476
rect 901 -1488 905 -1476
rect 827 -1493 855 -1488
rect 863 -1493 893 -1488
rect 901 -1493 915 -1488
rect 804 -1501 824 -1496
rect 827 -1501 831 -1493
rect 863 -1496 867 -1493
rect 901 -1496 905 -1493
rect 342 -1512 412 -1509
rect 342 -1516 345 -1512
rect 349 -1516 405 -1512
rect 409 -1516 412 -1512
rect 342 -1518 412 -1516
rect 352 -1524 356 -1518
rect 390 -1524 394 -1518
rect 288 -1551 316 -1546
rect 316 -1576 320 -1574
rect 270 -1581 320 -1576
rect 809 -1533 819 -1528
rect 855 -1530 859 -1516
rect 893 -1530 897 -1516
rect 845 -1532 915 -1530
rect 471 -1542 541 -1539
rect 471 -1546 474 -1542
rect 478 -1546 534 -1542
rect 538 -1546 541 -1542
rect 471 -1548 541 -1546
rect 324 -1576 328 -1574
rect 360 -1576 364 -1564
rect 398 -1576 402 -1564
rect 481 -1554 485 -1548
rect 519 -1554 523 -1548
rect 324 -1581 352 -1576
rect 360 -1581 390 -1576
rect 398 -1581 445 -1576
rect 324 -1589 328 -1581
rect 360 -1584 364 -1581
rect 398 -1584 402 -1581
rect 316 -1618 320 -1609
rect 352 -1618 356 -1604
rect 390 -1618 394 -1604
rect 445 -1606 449 -1604
rect 425 -1611 449 -1606
rect 453 -1606 457 -1604
rect 489 -1606 493 -1594
rect 527 -1606 531 -1594
rect 579 -1603 675 -1600
rect 453 -1611 481 -1606
rect 489 -1611 519 -1606
rect 527 -1611 574 -1606
rect 306 -1620 412 -1618
rect 306 -1624 308 -1620
rect 312 -1624 406 -1620
rect 410 -1624 412 -1620
rect 306 -1626 412 -1624
rect 425 -1641 431 -1611
rect 453 -1619 457 -1611
rect 489 -1614 493 -1611
rect 527 -1614 531 -1611
rect 261 -1646 431 -1641
rect 445 -1648 449 -1639
rect 481 -1648 485 -1634
rect 519 -1648 523 -1634
rect 435 -1650 541 -1648
rect 435 -1654 437 -1650
rect 441 -1654 535 -1650
rect 539 -1654 541 -1650
rect 435 -1656 541 -1654
rect 569 -1675 574 -1611
rect 579 -1607 608 -1603
rect 612 -1607 668 -1603
rect 672 -1607 675 -1603
rect 579 -1609 675 -1607
rect 579 -1645 583 -1609
rect 615 -1615 619 -1609
rect 653 -1615 657 -1609
rect 587 -1667 591 -1665
rect 623 -1667 627 -1655
rect 661 -1667 665 -1655
rect 587 -1672 615 -1667
rect 623 -1672 653 -1667
rect 661 -1672 698 -1667
rect 345 -1682 415 -1679
rect 569 -1680 584 -1675
rect 587 -1680 591 -1672
rect 623 -1675 627 -1672
rect 661 -1675 665 -1672
rect 345 -1686 348 -1682
rect 352 -1686 408 -1682
rect 412 -1686 415 -1682
rect 345 -1688 415 -1686
rect 355 -1694 359 -1688
rect 393 -1694 397 -1688
rect 288 -1721 319 -1716
rect 319 -1746 323 -1744
rect 270 -1751 323 -1746
rect 476 -1712 546 -1709
rect 476 -1716 479 -1712
rect 483 -1716 539 -1712
rect 543 -1716 546 -1712
rect 476 -1718 546 -1716
rect 569 -1712 579 -1707
rect 615 -1709 619 -1695
rect 653 -1709 657 -1695
rect 605 -1711 675 -1709
rect 327 -1746 331 -1744
rect 363 -1746 367 -1734
rect 401 -1746 405 -1734
rect 486 -1724 490 -1718
rect 524 -1724 528 -1718
rect 327 -1751 355 -1746
rect 363 -1751 393 -1746
rect 401 -1751 450 -1746
rect 327 -1759 331 -1751
rect 363 -1754 367 -1751
rect 401 -1754 405 -1751
rect 319 -1788 323 -1779
rect 355 -1788 359 -1774
rect 393 -1788 397 -1774
rect 450 -1776 454 -1774
rect 420 -1781 454 -1776
rect 458 -1776 462 -1774
rect 494 -1776 498 -1764
rect 532 -1776 536 -1764
rect 569 -1776 574 -1712
rect 605 -1715 607 -1711
rect 611 -1715 669 -1711
rect 673 -1715 675 -1711
rect 605 -1717 675 -1715
rect 458 -1781 486 -1776
rect 494 -1781 524 -1776
rect 532 -1781 574 -1776
rect 309 -1790 415 -1788
rect 309 -1794 311 -1790
rect 315 -1794 409 -1790
rect 413 -1794 415 -1790
rect 309 -1796 415 -1794
rect 345 -1826 415 -1823
rect 345 -1830 348 -1826
rect 352 -1830 408 -1826
rect 412 -1830 415 -1826
rect 345 -1832 415 -1830
rect 355 -1838 359 -1832
rect 393 -1838 397 -1832
rect 252 -1865 319 -1860
rect 319 -1890 323 -1888
rect 243 -1895 323 -1890
rect 327 -1890 331 -1888
rect 363 -1890 367 -1878
rect 401 -1890 405 -1878
rect 420 -1890 425 -1781
rect 458 -1789 462 -1781
rect 494 -1784 498 -1781
rect 532 -1784 536 -1781
rect 450 -1818 454 -1809
rect 486 -1818 490 -1804
rect 524 -1818 528 -1804
rect 440 -1820 546 -1818
rect 440 -1824 442 -1820
rect 446 -1824 540 -1820
rect 544 -1824 546 -1820
rect 440 -1826 546 -1824
rect 693 -1864 698 -1672
rect 708 -1792 804 -1789
rect 708 -1796 737 -1792
rect 741 -1796 797 -1792
rect 801 -1796 804 -1792
rect 708 -1798 804 -1796
rect 708 -1834 712 -1798
rect 744 -1804 748 -1798
rect 782 -1804 786 -1798
rect 716 -1856 720 -1854
rect 752 -1856 756 -1844
rect 790 -1856 794 -1844
rect 809 -1856 814 -1533
rect 845 -1536 847 -1532
rect 851 -1536 909 -1532
rect 913 -1536 915 -1532
rect 845 -1538 915 -1536
rect 716 -1861 744 -1856
rect 752 -1861 782 -1856
rect 790 -1861 814 -1856
rect 693 -1869 713 -1864
rect 716 -1869 720 -1861
rect 752 -1864 756 -1861
rect 790 -1864 794 -1861
rect 327 -1895 355 -1890
rect 363 -1895 393 -1890
rect 401 -1895 425 -1890
rect 327 -1903 331 -1895
rect 363 -1898 367 -1895
rect 401 -1898 405 -1895
rect 693 -1901 708 -1896
rect 744 -1898 748 -1884
rect 782 -1898 786 -1884
rect 734 -1900 804 -1898
rect 319 -1932 323 -1923
rect 355 -1932 359 -1918
rect 393 -1932 397 -1918
rect 309 -1934 415 -1932
rect 309 -1938 311 -1934
rect 315 -1938 409 -1934
rect 413 -1938 415 -1934
rect 309 -1940 415 -1938
rect 345 -1953 415 -1950
rect 345 -1957 348 -1953
rect 352 -1957 408 -1953
rect 412 -1957 415 -1953
rect 345 -1959 415 -1957
rect 355 -1965 359 -1959
rect 393 -1965 397 -1959
rect 288 -1992 319 -1987
rect 319 -2017 323 -2015
rect 270 -2022 323 -2017
rect 476 -1983 546 -1980
rect 476 -1987 479 -1983
rect 483 -1987 539 -1983
rect 543 -1987 546 -1983
rect 476 -1989 546 -1987
rect 327 -2017 331 -2015
rect 363 -2017 367 -2005
rect 401 -2017 405 -2005
rect 486 -1995 490 -1989
rect 524 -1995 528 -1989
rect 327 -2022 355 -2017
rect 363 -2022 393 -2017
rect 401 -2022 450 -2017
rect 327 -2030 331 -2022
rect 363 -2025 367 -2022
rect 401 -2025 405 -2022
rect 319 -2059 323 -2050
rect 355 -2059 359 -2045
rect 393 -2059 397 -2045
rect 450 -2047 454 -2045
rect 420 -2052 454 -2047
rect 611 -2013 681 -2010
rect 611 -2017 614 -2013
rect 618 -2017 674 -2013
rect 678 -2017 681 -2013
rect 611 -2019 681 -2017
rect 458 -2047 462 -2045
rect 494 -2047 498 -2035
rect 532 -2047 536 -2035
rect 621 -2025 625 -2019
rect 659 -2025 663 -2019
rect 458 -2052 486 -2047
rect 494 -2052 524 -2047
rect 532 -2052 585 -2047
rect 309 -2061 415 -2059
rect 309 -2065 311 -2061
rect 315 -2065 409 -2061
rect 413 -2065 415 -2061
rect 309 -2067 415 -2065
rect 345 -2097 415 -2094
rect 345 -2101 348 -2097
rect 352 -2101 408 -2097
rect 412 -2101 415 -2097
rect 345 -2103 415 -2101
rect 355 -2109 359 -2103
rect 393 -2109 397 -2103
rect 252 -2136 319 -2131
rect 319 -2161 323 -2159
rect 234 -2166 323 -2161
rect 327 -2161 331 -2159
rect 363 -2161 367 -2149
rect 401 -2161 405 -2149
rect 420 -2161 425 -2052
rect 458 -2060 462 -2052
rect 494 -2055 498 -2052
rect 532 -2055 536 -2052
rect 450 -2089 454 -2080
rect 486 -2089 490 -2075
rect 524 -2089 528 -2075
rect 585 -2077 589 -2075
rect 558 -2082 589 -2077
rect 593 -2077 597 -2075
rect 629 -2077 633 -2065
rect 667 -2077 671 -2065
rect 693 -2077 698 -1901
rect 734 -1904 736 -1900
rect 740 -1904 798 -1900
rect 802 -1904 804 -1900
rect 734 -1906 804 -1904
rect 593 -2082 621 -2077
rect 629 -2082 659 -2077
rect 667 -2082 698 -2077
rect 440 -2091 546 -2089
rect 440 -2095 442 -2091
rect 446 -2095 540 -2091
rect 544 -2095 546 -2091
rect 440 -2097 546 -2095
rect 327 -2166 355 -2161
rect 363 -2166 393 -2161
rect 401 -2166 425 -2161
rect 327 -2174 331 -2166
rect 363 -2169 367 -2166
rect 401 -2169 405 -2166
rect 319 -2203 323 -2194
rect 355 -2203 359 -2189
rect 393 -2203 397 -2189
rect 309 -2205 415 -2203
rect 309 -2209 311 -2205
rect 315 -2209 409 -2205
rect 413 -2209 415 -2205
rect 309 -2211 415 -2209
rect 558 -2220 563 -2082
rect 593 -2090 597 -2082
rect 629 -2085 633 -2082
rect 667 -2085 671 -2082
rect 585 -2119 589 -2110
rect 621 -2119 625 -2105
rect 659 -2119 663 -2105
rect 575 -2121 681 -2119
rect 575 -2125 577 -2121
rect 581 -2125 675 -2121
rect 679 -2125 681 -2121
rect 575 -2127 681 -2125
rect 225 -2225 563 -2220
<< m2contact >>
rect 220 280 225 285
rect 229 230 234 235
rect 58 95 63 100
rect 90 95 95 100
rect 238 91 243 96
rect 229 1 234 6
rect 220 -29 225 -24
rect 489 49 494 54
rect 247 -86 252 -81
rect 464 -86 469 -81
rect 58 -195 63 -190
rect 90 -195 95 -190
rect 256 -199 261 -194
rect 238 -289 243 -284
rect 247 -319 252 -314
rect 220 -415 225 -410
rect 229 -445 234 -440
rect 691 -363 696 -358
rect 247 -511 252 -505
rect 265 -533 270 -528
rect 645 -533 650 -528
rect 58 -612 63 -607
rect 90 -612 95 -607
rect 274 -616 279 -611
rect 256 -706 261 -701
rect 265 -736 270 -731
rect 238 -850 243 -845
rect 247 -880 252 -875
rect 265 -945 270 -940
rect 890 -795 895 -790
rect 220 -1020 225 -1015
rect 229 -1050 234 -1045
rect 247 -1164 252 -1159
rect 265 -1194 270 -1189
rect 283 -1249 288 -1244
rect 853 -1249 858 -1244
rect 58 -1313 63 -1308
rect 90 -1313 95 -1308
rect 274 -1407 279 -1402
rect 283 -1437 288 -1432
rect 283 -1551 288 -1546
rect 265 -1581 270 -1576
rect 256 -1646 261 -1641
rect 283 -1721 288 -1716
rect 265 -1751 270 -1746
rect 247 -1865 252 -1860
rect 238 -1895 243 -1890
rect 283 -1992 288 -1987
rect 265 -2022 270 -2017
rect 247 -2136 252 -2131
rect 229 -2166 234 -2161
rect 220 -2225 225 -2220
<< metal2 >>
rect 63 95 90 100
rect 220 -24 225 280
rect 63 -195 90 -190
rect 220 -410 225 -29
rect 63 -612 90 -607
rect 220 -1015 225 -415
rect 63 -1313 90 -1308
rect 220 -2220 225 -1020
rect 229 6 234 230
rect 229 -440 234 1
rect 229 -1045 234 -445
rect 229 -2161 234 -1050
rect 238 -284 243 91
rect 464 49 489 54
rect 464 -81 469 49
rect 238 -845 243 -289
rect 238 -1890 243 -850
rect 247 -314 252 -86
rect 247 -505 252 -319
rect 247 -875 252 -511
rect 247 -1159 252 -880
rect 247 -1860 252 -1164
rect 256 -701 261 -199
rect 645 -363 691 -358
rect 645 -528 650 -363
rect 256 -1641 261 -706
rect 265 -731 270 -533
rect 265 -940 270 -736
rect 265 -1189 270 -945
rect 265 -1576 270 -1194
rect 274 -1402 279 -616
rect 853 -795 890 -790
rect 853 -1244 858 -795
rect 247 -2131 252 -1865
rect 265 -1746 270 -1581
rect 265 -2017 270 -1751
rect 283 -1432 288 -1249
rect 283 -1546 288 -1437
rect 283 -1716 288 -1551
rect 283 -1987 288 -1721
<< labels >>
rlabel metal1 -5 -35 -5 -35 3 vdd
rlabel metal1 97 -34 97 -34 7 gnd
rlabel metal1 97 17 97 17 7 gnd
rlabel metal1 -5 16 -5 16 3 vdd
rlabel metal1 149 39 149 39 5 vdd
rlabel metal1 149 159 149 159 5 vdd
rlabel metal1 148 57 148 57 1 gnd
rlabel metal1 187 159 187 159 5 vdd
rlabel metal1 186 57 186 57 1 gnd
rlabel metal1 111 64 111 64 1 gnd
rlabel metal1 148 -63 148 -63 1 gnd
rlabel metal1 88 -13 88 -13 1 b0
rlabel metal1 60 0 60 0 1 a0_not
rlabel metal1 85 -59 85 -59 1 b0_not
rlabel metal1 60 25 60 25 1 a0
rlabel metal1 130 -13 130 -13 1 p0_not
rlabel metal1 160 -26 160 -26 1 p0
rlabel metal1 135 94 135 94 1 g0_mid
rlabel metal1 169 94 169 94 1 g0_not
rlabel metal1 200 94 200 94 1 g0
rlabel metal1 -5 -325 -5 -325 3 vdd
rlabel metal1 97 -324 97 -324 7 gnd
rlabel metal1 97 -273 97 -273 7 gnd
rlabel metal1 -5 -274 -5 -274 3 vdd
rlabel metal1 149 -251 149 -251 5 vdd
rlabel metal1 148 -353 148 -353 1 gnd
rlabel metal1 149 -131 149 -131 5 vdd
rlabel metal1 148 -233 148 -233 1 gnd
rlabel metal1 187 -131 187 -131 5 vdd
rlabel metal1 186 -233 186 -233 1 gnd
rlabel metal1 111 -226 111 -226 1 gnd
rlabel metal1 200 -196 200 -196 1 g1
rlabel metal1 169 -196 169 -196 1 g1_not
rlabel metal1 135 -196 135 -196 1 g1_mid
rlabel metal1 60 -265 60 -265 1 a1
rlabel metal1 60 -290 60 -290 1 a1_not
rlabel metal1 88 -303 88 -303 1 b1
rlabel metal1 85 -349 85 -349 1 b1_not
rlabel metal1 130 -303 130 -303 1 p1_not
rlabel metal1 160 -316 160 -316 1 p1
rlabel metal1 111 -643 111 -643 1 gnd
rlabel metal1 186 -650 186 -650 1 gnd
rlabel metal1 187 -548 187 -548 5 vdd
rlabel metal1 148 -650 148 -650 1 gnd
rlabel metal1 149 -548 149 -548 5 vdd
rlabel metal1 148 -770 148 -770 1 gnd
rlabel metal1 149 -668 149 -668 5 vdd
rlabel metal1 -5 -691 -5 -691 3 vdd
rlabel metal1 97 -690 97 -690 7 gnd
rlabel metal1 97 -741 97 -741 7 gnd
rlabel metal1 -5 -742 -5 -742 3 vdd
rlabel metal1 135 -613 135 -613 1 g2_mid
rlabel metal1 169 -613 169 -613 1 g2_not
rlabel metal1 200 -613 200 -613 1 g2
rlabel metal1 160 -733 160 -733 1 p2
rlabel metal1 130 -720 130 -720 1 p2_not
rlabel metal1 60 -682 60 -682 1 a2
rlabel metal1 60 -707 60 -707 1 a2_not
rlabel metal1 85 -766 85 -766 1 b2_not
rlabel metal1 88 -720 88 -720 1 b2
rlabel metal1 365 -27 365 -27 1 w1
rlabel metal1 333 38 333 38 5 vdd
rlabel metal1 318 -70 318 -70 1 gnd
rlabel metal1 257 210 257 210 3 vdd
rlabel metal1 359 211 359 211 7 gnd
rlabel metal1 359 262 359 262 7 gnd
rlabel metal1 257 261 257 261 3 vdd
rlabel metal1 411 284 411 284 5 vdd
rlabel metal1 410 182 410 182 1 gnd
rlabel metal1 423 218 423 218 7 s0
rlabel metal1 424 58 424 58 1 gnd
rlabel metal1 439 166 439 166 5 vdd
rlabel metal1 473 101 473 101 1 c1
rlabel metal1 493 29 493 29 3 vdd
rlabel metal1 595 30 595 30 7 gnd
rlabel metal1 595 81 595 81 7 gnd
rlabel metal1 493 80 493 80 3 vdd
rlabel metal1 647 103 647 103 5 vdd
rlabel metal1 646 1 646 1 1 gnd
rlabel metal1 660 38 660 38 7 s1
rlabel metal1 413 -252 413 -252 5 vdd
rlabel metal1 398 -360 398 -360 1 gnd
rlabel metal1 255 -27 255 -27 1 p0
rlabel metal1 249 3 249 3 1 c0
rlabel metal1 328 -286 328 -286 1 g0
rlabel metal1 328 -317 328 -317 1 p1
rlabel metal1 326 -486 326 -486 1 gnd
rlabel metal1 341 -378 341 -378 5 vdd
rlabel metal1 270 -413 270 -413 1 p0
rlabel metal1 270 -443 270 -443 1 c0
rlabel metal1 455 -516 455 -516 1 gnd
rlabel metal1 470 -408 470 -408 5 vdd
rlabel metal1 513 -473 513 -473 1 p1p0c0
rlabel metal1 457 -256 457 -256 1 p1g0
rlabel metal1 501 -232 501 -232 1 gnd
rlabel metal1 516 -124 516 -124 5 vdd
rlabel metal1 365 -669 365 -669 5 vdd
rlabel metal1 350 -777 350 -777 1 gnd
rlabel metal1 350 -921 350 -921 1 gnd
rlabel metal1 365 -813 365 -813 5 vdd
rlabel metal1 479 -951 479 -951 1 gnd
rlabel metal1 494 -843 494 -843 5 vdd
rlabel metal1 368 -983 368 -983 5 vdd
rlabel metal1 353 -1091 353 -1091 1 gnd
rlabel metal1 368 -1127 368 -1127 5 vdd
rlabel metal1 353 -1235 353 -1235 1 gnd
rlabel nwell 187 -1306 187 -1306 5 vdd
rlabel nwell 149 -1306 149 -1306 5 vdd
rlabel metal1 484 -1121 484 -1121 1 gnd
rlabel metal1 499 -1013 499 -1013 5 vdd
rlabel metal1 673 -541 673 -541 5 vdd
rlabel metal1 658 -649 658 -649 1 gnd
rlabel metal1 669 -897 669 -897 5 vdd
rlabel metal1 654 -1005 654 -1005 1 gnd
rlabel metal1 840 -678 840 -678 5 vdd
rlabel metal1 825 -786 825 -786 1 gnd
rlabel metal1 667 -310 667 -310 1 c2
rlabel metal1 621 -354 621 -354 1 gnd
rlabel metal1 636 -246 636 -246 5 vdd
rlabel metal1 695 -383 695 -383 3 vdd
rlabel metal1 797 -382 797 -382 7 gnd
rlabel metal1 797 -331 797 -331 7 gnd
rlabel metal1 695 -332 695 -332 3 vdd
rlabel metal1 849 -309 849 -309 5 vdd
rlabel metal1 848 -411 848 -411 1 gnd
rlabel metal1 863 -375 863 -375 7 s2
rlabel metal1 873 -743 873 -743 7 c3
rlabel metal1 1047 -843 1047 -843 1 gnd
rlabel metal1 1048 -741 1048 -741 5 vdd
rlabel metal1 894 -764 894 -764 3 vdd
rlabel metal1 996 -763 996 -763 7 gnd
rlabel metal1 996 -814 996 -814 7 gnd
rlabel metal1 894 -815 894 -815 3 vdd
rlabel metal1 1062 -807 1062 -807 7 s3
rlabel metal1 111 -1344 111 -1344 1 gnd
rlabel metal1 186 -1351 186 -1351 1 gnd
rlabel metal1 148 -1351 148 -1351 1 gnd
rlabel metal1 148 -1471 148 -1471 1 gnd
rlabel metal1 149 -1369 149 -1369 5 vdd
rlabel metal1 -5 -1392 -5 -1392 3 vdd
rlabel metal1 97 -1391 97 -1391 7 gnd
rlabel metal1 97 -1442 97 -1442 7 gnd
rlabel metal1 -5 -1443 -5 -1443 3 vdd
rlabel metal1 135 -1314 135 -1314 1 g3_mid
rlabel metal1 169 -1314 169 -1314 1 g3_not
rlabel metal1 200 -1314 200 -1314 1 g3
rlabel metal1 160 -1434 160 -1434 1 p3
rlabel metal1 60 -1383 60 -1383 1 a3
rlabel metal1 60 -1408 60 -1408 1 a3_not
rlabel metal1 85 -1467 85 -1467 1 b3_not
rlabel metal1 88 -1421 88 -1421 1 b3
rlabel metal1 130 -1421 130 -1421 1 p3_not
rlabel metal1 149 -1249 149 -1249 5 vdd
rlabel metal1 187 -1249 187 -1249 5 vdd
rlabel metal1 511 -1714 511 -1714 5 vdd
rlabel metal1 496 -1822 496 -1822 1 gnd
rlabel metal1 365 -1936 365 -1936 1 gnd
rlabel metal1 380 -1828 380 -1828 5 vdd
rlabel metal1 365 -1792 365 -1792 1 gnd
rlabel metal1 380 -1684 380 -1684 5 vdd
rlabel metal1 506 -1544 506 -1544 5 vdd
rlabel metal1 491 -1652 491 -1652 1 gnd
rlabel metal1 377 -1514 377 -1514 5 vdd
rlabel metal1 362 -1622 362 -1622 1 gnd
rlabel metal1 362 -1478 362 -1478 1 gnd
rlabel metal1 377 -1370 377 -1370 5 vdd
rlabel metal1 511 -1985 511 -1985 5 vdd
rlabel metal1 496 -2093 496 -2093 1 gnd
rlabel metal1 365 -2207 365 -2207 1 gnd
rlabel metal1 380 -2099 380 -2099 5 vdd
rlabel metal1 365 -2063 365 -2063 1 gnd
rlabel metal1 380 -1955 380 -1955 5 vdd
rlabel metal1 646 -2015 646 -2015 5 vdd
rlabel metal1 631 -2123 631 -2123 1 gnd
rlabel metal1 516 -1438 516 -1438 1 gnd
rlabel metal1 531 -1330 531 -1330 5 vdd
rlabel metal1 640 -1605 640 -1605 5 vdd
rlabel metal1 625 -1713 625 -1713 1 gnd
rlabel metal1 769 -1794 769 -1794 5 vdd
rlabel metal1 754 -1902 754 -1902 1 gnd
rlabel metal1 865 -1534 865 -1534 1 gnd
rlabel metal1 880 -1426 880 -1426 5 vdd
rlabel metal1 912 -1491 912 -1491 1 cout
<< end >>
