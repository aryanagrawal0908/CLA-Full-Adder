magic
tech scmos
timestamp 1732033240
<< nwell >>
rect -354 117 -322 243
rect -302 117 -270 243
rect -250 179 -218 243
rect -198 179 -166 243
rect -153 187 -89 251
rect 889 245 953 277
rect 889 194 953 226
rect 1031 224 1063 288
rect 1132 225 1164 351
rect 1184 225 1216 351
rect 1236 287 1268 351
rect 1288 287 1320 351
rect 1333 295 1397 359
rect 1403 295 1435 339
rect 133 99 165 163
rect 171 99 203 163
rect 404 107 474 171
rect 368 64 400 98
rect 889 64 953 96
rect -355 -94 -323 32
rect -303 -94 -271 32
rect -251 -32 -219 32
rect -199 -32 -167 32
rect -154 -24 -90 40
rect -9 0 55 32
rect -9 -51 55 -19
rect 133 -21 165 43
rect 298 -21 368 43
rect 889 13 953 45
rect 1031 43 1063 107
rect 1131 25 1163 151
rect 1183 25 1215 151
rect 1235 87 1267 151
rect 1287 87 1319 151
rect 1332 95 1396 159
rect 1402 95 1434 139
rect 262 -64 294 -30
rect -363 -298 -331 -172
rect -311 -298 -279 -172
rect -259 -236 -227 -172
rect -207 -236 -175 -172
rect -162 -228 -98 -164
rect 133 -191 165 -127
rect 171 -191 203 -127
rect 481 -183 551 -119
rect 445 -226 477 -192
rect -9 -290 55 -258
rect -9 -341 55 -309
rect 133 -311 165 -247
rect 378 -311 448 -247
rect 601 -305 671 -241
rect 342 -354 374 -320
rect 565 -348 597 -314
rect 889 -348 953 -316
rect -364 -509 -332 -383
rect -312 -509 -280 -383
rect -260 -447 -228 -383
rect -208 -447 -176 -383
rect -163 -439 -99 -375
rect 306 -437 376 -373
rect 889 -399 953 -367
rect 1031 -369 1063 -305
rect 1130 -374 1162 -248
rect 1182 -374 1214 -248
rect 1234 -312 1266 -248
rect 1286 -312 1318 -248
rect 1331 -304 1395 -240
rect 1401 -304 1433 -260
rect 270 -480 302 -446
rect 435 -467 505 -403
rect 399 -510 431 -476
rect -369 -704 -337 -578
rect -317 -704 -285 -578
rect -265 -642 -233 -578
rect -213 -642 -181 -578
rect -168 -634 -104 -570
rect 133 -608 165 -544
rect 171 -608 203 -544
rect 638 -600 708 -536
rect 602 -643 634 -609
rect -9 -707 55 -675
rect -9 -758 55 -726
rect 133 -728 165 -664
rect 330 -728 400 -664
rect 805 -737 875 -673
rect 294 -771 326 -737
rect 769 -780 801 -746
rect 890 -780 954 -748
rect -370 -915 -338 -789
rect -318 -915 -286 -789
rect -266 -853 -234 -789
rect -214 -853 -182 -789
rect -169 -845 -105 -781
rect 330 -872 400 -808
rect 890 -831 954 -799
rect 1032 -801 1064 -737
rect 1130 -788 1162 -662
rect 1182 -788 1214 -662
rect 1234 -726 1266 -662
rect 1286 -726 1318 -662
rect 1331 -718 1395 -654
rect 1401 -718 1433 -674
rect 294 -915 326 -881
rect 459 -902 529 -838
rect 423 -945 455 -911
rect 634 -956 704 -892
rect 333 -1042 403 -978
rect 598 -999 630 -965
rect 297 -1085 329 -1051
rect 464 -1072 534 -1008
rect 428 -1115 460 -1081
rect 333 -1186 403 -1122
rect 297 -1229 329 -1195
rect -356 -1406 -324 -1280
rect -304 -1406 -272 -1280
rect -252 -1344 -220 -1280
rect -200 -1344 -168 -1280
rect -155 -1336 -91 -1272
rect 133 -1309 165 -1245
rect 171 -1309 203 -1245
rect -9 -1408 55 -1376
rect -9 -1459 55 -1427
rect 133 -1429 165 -1365
rect 342 -1429 412 -1365
rect 496 -1389 566 -1325
rect 460 -1432 492 -1398
rect 306 -1472 338 -1438
rect -357 -1617 -325 -1491
rect -305 -1617 -273 -1491
rect -253 -1555 -221 -1491
rect -201 -1555 -169 -1491
rect -156 -1547 -92 -1483
rect 845 -1485 915 -1421
rect 1131 -1484 1163 -1358
rect 1183 -1484 1215 -1358
rect 1235 -1422 1267 -1358
rect 1287 -1422 1319 -1358
rect 1332 -1414 1396 -1350
rect 1402 -1414 1434 -1370
rect 342 -1573 412 -1509
rect 809 -1528 841 -1494
rect 306 -1616 338 -1582
rect 471 -1603 541 -1539
rect 435 -1646 467 -1612
rect 605 -1664 675 -1600
rect 345 -1743 415 -1679
rect 569 -1707 601 -1673
rect 309 -1786 341 -1752
rect 476 -1773 546 -1709
rect 440 -1816 472 -1782
rect 345 -1887 415 -1823
rect 734 -1853 804 -1789
rect 698 -1896 730 -1862
rect 309 -1930 341 -1896
rect 345 -2014 415 -1950
rect 309 -2057 341 -2023
rect 476 -2044 546 -1980
rect 440 -2087 472 -2053
rect 611 -2074 681 -2010
rect 345 -2158 415 -2094
rect 575 -2117 607 -2083
rect 309 -2201 341 -2167
<< ntransistor >>
rect 964 260 984 262
rect 1014 252 1016 272
rect 1014 220 1016 240
rect 1348 264 1350 284
rect 1380 264 1382 284
rect 1418 274 1420 284
rect 1251 240 1253 260
rect 1303 240 1305 260
rect 964 209 984 211
rect 1046 193 1048 213
rect 1147 193 1149 213
rect 1199 193 1201 213
rect 1251 193 1253 213
rect 1303 193 1305 213
rect -138 156 -136 176
rect -106 156 -104 176
rect -235 132 -233 152
rect -183 132 -181 152
rect -339 85 -337 105
rect -287 85 -285 105
rect -235 85 -233 105
rect -183 85 -181 105
rect 116 101 118 121
rect 116 69 118 89
rect 383 106 385 126
rect 148 68 150 88
rect 186 68 188 88
rect 419 76 421 96
rect 457 76 459 96
rect 964 79 984 81
rect 1014 71 1016 91
rect 1014 39 1016 59
rect 1347 64 1349 84
rect 1379 64 1381 84
rect 1417 74 1419 84
rect 1250 40 1252 60
rect 1302 40 1304 60
rect 964 28 984 30
rect 66 15 86 17
rect 116 7 118 27
rect 116 -25 118 -5
rect 277 -22 279 -2
rect 1046 12 1048 32
rect 1146 -7 1148 13
rect 1198 -7 1200 13
rect 1250 -7 1252 13
rect 1302 -7 1304 13
rect -139 -55 -137 -35
rect -107 -55 -105 -35
rect 66 -36 86 -34
rect 148 -52 150 -32
rect 313 -52 315 -32
rect 351 -52 353 -32
rect -236 -79 -234 -59
rect -184 -79 -182 -59
rect -340 -126 -338 -106
rect -288 -126 -286 -106
rect -236 -126 -234 -106
rect -184 -126 -182 -106
rect 116 -189 118 -169
rect 116 -221 118 -201
rect 460 -184 462 -164
rect 148 -222 150 -202
rect 186 -222 188 -202
rect 496 -214 498 -194
rect 534 -214 536 -194
rect -147 -259 -145 -239
rect -115 -259 -113 -239
rect -244 -283 -242 -263
rect -192 -283 -190 -263
rect 66 -275 86 -273
rect 116 -283 118 -263
rect -348 -330 -346 -310
rect -296 -330 -294 -310
rect -244 -330 -242 -310
rect -192 -330 -190 -310
rect 116 -315 118 -295
rect 357 -312 359 -292
rect 66 -326 86 -324
rect 148 -342 150 -322
rect 580 -306 582 -286
rect 393 -342 395 -322
rect 431 -342 433 -322
rect 616 -336 618 -316
rect 654 -336 656 -316
rect 964 -333 984 -331
rect 1014 -341 1016 -321
rect 1014 -373 1016 -353
rect 1346 -335 1348 -315
rect 1378 -335 1380 -315
rect 1416 -325 1418 -315
rect 1249 -359 1251 -339
rect 1301 -359 1303 -339
rect 964 -384 984 -382
rect 285 -438 287 -418
rect 1046 -400 1048 -380
rect 1145 -406 1147 -386
rect 1197 -406 1199 -386
rect 1249 -406 1251 -386
rect 1301 -406 1303 -386
rect -148 -470 -146 -450
rect -116 -470 -114 -450
rect 321 -468 323 -448
rect 359 -468 361 -448
rect 414 -468 416 -448
rect -245 -494 -243 -474
rect -193 -494 -191 -474
rect 450 -498 452 -478
rect 488 -498 490 -478
rect -349 -541 -347 -521
rect -297 -541 -295 -521
rect -245 -541 -243 -521
rect -193 -541 -191 -521
rect 116 -606 118 -586
rect 116 -638 118 -618
rect 617 -601 619 -581
rect -153 -665 -151 -645
rect -121 -665 -119 -645
rect 148 -639 150 -619
rect 186 -639 188 -619
rect 653 -631 655 -611
rect 691 -631 693 -611
rect -250 -689 -248 -669
rect -198 -689 -196 -669
rect 66 -692 86 -690
rect 116 -700 118 -680
rect -354 -736 -352 -716
rect -302 -736 -300 -716
rect -250 -736 -248 -716
rect -198 -736 -196 -716
rect 116 -732 118 -712
rect 309 -729 311 -709
rect 66 -743 86 -741
rect 148 -759 150 -739
rect 784 -738 786 -718
rect 345 -759 347 -739
rect 383 -759 385 -739
rect 820 -768 822 -748
rect 858 -768 860 -748
rect 965 -765 985 -763
rect 1015 -773 1017 -753
rect 1015 -805 1017 -785
rect 1346 -749 1348 -729
rect 1378 -749 1380 -729
rect 1416 -739 1418 -729
rect 1249 -773 1251 -753
rect 1301 -773 1303 -753
rect 965 -816 985 -814
rect -154 -876 -152 -856
rect -122 -876 -120 -856
rect 309 -873 311 -853
rect 1047 -832 1049 -812
rect 1145 -820 1147 -800
rect 1197 -820 1199 -800
rect 1249 -820 1251 -800
rect 1301 -820 1303 -800
rect -251 -900 -249 -880
rect -199 -900 -197 -880
rect 345 -903 347 -883
rect 383 -903 385 -883
rect 438 -903 440 -883
rect -355 -947 -353 -927
rect -303 -947 -301 -927
rect -251 -947 -249 -927
rect -199 -947 -197 -927
rect 474 -933 476 -913
rect 512 -933 514 -913
rect 613 -957 615 -937
rect 649 -987 651 -967
rect 687 -987 689 -967
rect 312 -1043 314 -1023
rect 348 -1073 350 -1053
rect 386 -1073 388 -1053
rect 443 -1073 445 -1053
rect 479 -1103 481 -1083
rect 517 -1103 519 -1083
rect 312 -1187 314 -1167
rect 348 -1217 350 -1197
rect 386 -1217 388 -1197
rect 116 -1307 118 -1287
rect 116 -1339 118 -1319
rect -140 -1367 -138 -1347
rect -108 -1367 -106 -1347
rect 148 -1340 150 -1320
rect 186 -1340 188 -1320
rect -237 -1391 -235 -1371
rect -185 -1391 -183 -1371
rect 66 -1393 86 -1391
rect 116 -1401 118 -1381
rect -341 -1438 -339 -1418
rect -289 -1438 -287 -1418
rect -237 -1438 -235 -1418
rect -185 -1438 -183 -1418
rect 116 -1433 118 -1413
rect 321 -1430 323 -1410
rect 475 -1390 477 -1370
rect 66 -1444 86 -1442
rect 148 -1460 150 -1440
rect 511 -1420 513 -1400
rect 549 -1420 551 -1400
rect 357 -1460 359 -1440
rect 395 -1460 397 -1440
rect 824 -1486 826 -1466
rect 1347 -1445 1349 -1425
rect 1379 -1445 1381 -1425
rect 1417 -1435 1419 -1425
rect 1250 -1469 1252 -1449
rect 1302 -1469 1304 -1449
rect 860 -1516 862 -1496
rect 898 -1516 900 -1496
rect 1146 -1516 1148 -1496
rect 1198 -1516 1200 -1496
rect 1250 -1516 1252 -1496
rect 1302 -1516 1304 -1496
rect -141 -1578 -139 -1558
rect -109 -1578 -107 -1558
rect 321 -1574 323 -1554
rect -238 -1602 -236 -1582
rect -186 -1602 -184 -1582
rect 357 -1604 359 -1584
rect 395 -1604 397 -1584
rect 450 -1604 452 -1584
rect -342 -1649 -340 -1629
rect -290 -1649 -288 -1629
rect -238 -1649 -236 -1629
rect -186 -1649 -184 -1629
rect 486 -1634 488 -1614
rect 524 -1634 526 -1614
rect 584 -1665 586 -1645
rect 324 -1744 326 -1724
rect 620 -1695 622 -1675
rect 658 -1695 660 -1675
rect 360 -1774 362 -1754
rect 398 -1774 400 -1754
rect 455 -1774 457 -1754
rect 491 -1804 493 -1784
rect 529 -1804 531 -1784
rect 324 -1888 326 -1868
rect 713 -1854 715 -1834
rect 749 -1884 751 -1864
rect 787 -1884 789 -1864
rect 360 -1918 362 -1898
rect 398 -1918 400 -1898
rect 324 -2015 326 -1995
rect 360 -2045 362 -2025
rect 398 -2045 400 -2025
rect 455 -2045 457 -2025
rect 491 -2075 493 -2055
rect 529 -2075 531 -2055
rect 590 -2075 592 -2055
rect 324 -2159 326 -2139
rect 626 -2105 628 -2085
rect 664 -2105 666 -2085
rect 360 -2189 362 -2169
rect 398 -2189 400 -2169
<< ptransistor >>
rect 1147 296 1149 336
rect 1199 296 1201 336
rect 1251 296 1253 336
rect 1303 296 1305 336
rect 1348 304 1350 344
rect 1380 304 1382 344
rect 1418 304 1420 324
rect 904 260 944 262
rect -339 188 -337 228
rect -287 188 -285 228
rect -235 188 -233 228
rect -183 188 -181 228
rect -138 196 -136 236
rect -106 196 -104 236
rect 1046 233 1048 273
rect 1147 234 1149 274
rect 1199 234 1201 274
rect 904 209 944 211
rect -339 126 -337 166
rect -287 126 -285 166
rect 148 108 150 148
rect 186 108 188 148
rect 419 116 421 156
rect 457 116 459 156
rect 383 71 385 91
rect 1146 96 1148 136
rect 1198 96 1200 136
rect 1250 96 1252 136
rect 1302 96 1304 136
rect 1347 104 1349 144
rect 1379 104 1381 144
rect 1417 104 1419 124
rect 904 79 944 81
rect 1046 52 1048 92
rect 1146 34 1148 74
rect 1198 34 1200 74
rect 904 28 944 30
rect -340 -23 -338 17
rect -288 -23 -286 17
rect -236 -23 -234 17
rect -184 -23 -182 17
rect -139 -15 -137 25
rect -107 -15 -105 25
rect 6 15 46 17
rect 148 -12 150 28
rect 313 -12 315 28
rect 351 -12 353 28
rect -340 -85 -338 -45
rect -288 -85 -286 -45
rect 6 -36 46 -34
rect 277 -57 279 -37
rect -348 -227 -346 -187
rect -296 -227 -294 -187
rect -244 -227 -242 -187
rect -192 -227 -190 -187
rect -147 -219 -145 -179
rect -115 -219 -113 -179
rect 148 -182 150 -142
rect 186 -182 188 -142
rect 496 -174 498 -134
rect 534 -174 536 -134
rect 460 -219 462 -199
rect -348 -289 -346 -249
rect -296 -289 -294 -249
rect 6 -275 46 -273
rect 148 -302 150 -262
rect 393 -302 395 -262
rect 431 -302 433 -262
rect 6 -326 46 -324
rect 616 -296 618 -256
rect 654 -296 656 -256
rect 1145 -303 1147 -263
rect 1197 -303 1199 -263
rect 1249 -303 1251 -263
rect 1301 -303 1303 -263
rect 1346 -295 1348 -255
rect 1378 -295 1380 -255
rect 1416 -295 1418 -275
rect 357 -347 359 -327
rect 580 -341 582 -321
rect 904 -333 944 -331
rect 1046 -360 1048 -320
rect 1145 -365 1147 -325
rect 1197 -365 1199 -325
rect 904 -384 944 -382
rect -349 -438 -347 -398
rect -297 -438 -295 -398
rect -245 -438 -243 -398
rect -193 -438 -191 -398
rect -148 -430 -146 -390
rect -116 -430 -114 -390
rect 321 -428 323 -388
rect 359 -428 361 -388
rect -349 -500 -347 -460
rect -297 -500 -295 -460
rect 285 -473 287 -453
rect 450 -458 452 -418
rect 488 -458 490 -418
rect 414 -503 416 -483
rect -354 -633 -352 -593
rect -302 -633 -300 -593
rect -250 -633 -248 -593
rect -198 -633 -196 -593
rect -153 -625 -151 -585
rect -121 -625 -119 -585
rect 148 -599 150 -559
rect 186 -599 188 -559
rect 653 -591 655 -551
rect 691 -591 693 -551
rect -354 -695 -352 -655
rect -302 -695 -300 -655
rect 617 -636 619 -616
rect 6 -692 46 -690
rect 148 -719 150 -679
rect 345 -719 347 -679
rect 383 -719 385 -679
rect 6 -743 46 -741
rect 820 -728 822 -688
rect 858 -728 860 -688
rect 1145 -717 1147 -677
rect 1197 -717 1199 -677
rect 1249 -717 1251 -677
rect 1301 -717 1303 -677
rect 1346 -709 1348 -669
rect 1378 -709 1380 -669
rect 1416 -709 1418 -689
rect 309 -764 311 -744
rect 784 -773 786 -753
rect 905 -765 945 -763
rect -355 -844 -353 -804
rect -303 -844 -301 -804
rect -251 -844 -249 -804
rect -199 -844 -197 -804
rect -154 -836 -152 -796
rect -122 -836 -120 -796
rect 1047 -792 1049 -752
rect 1145 -779 1147 -739
rect 1197 -779 1199 -739
rect 905 -816 945 -814
rect -355 -906 -353 -866
rect -303 -906 -301 -866
rect 345 -863 347 -823
rect 383 -863 385 -823
rect 309 -908 311 -888
rect 474 -893 476 -853
rect 512 -893 514 -853
rect 438 -938 440 -918
rect 649 -947 651 -907
rect 687 -947 689 -907
rect 613 -992 615 -972
rect 348 -1033 350 -993
rect 386 -1033 388 -993
rect 312 -1078 314 -1058
rect 479 -1063 481 -1023
rect 517 -1063 519 -1023
rect 443 -1108 445 -1088
rect 348 -1177 350 -1137
rect 386 -1177 388 -1137
rect 312 -1222 314 -1202
rect -341 -1335 -339 -1295
rect -289 -1335 -287 -1295
rect -237 -1335 -235 -1295
rect -185 -1335 -183 -1295
rect -140 -1327 -138 -1287
rect -108 -1327 -106 -1287
rect 148 -1300 150 -1260
rect 186 -1300 188 -1260
rect -341 -1397 -339 -1357
rect -289 -1397 -287 -1357
rect 6 -1393 46 -1391
rect 148 -1420 150 -1380
rect 357 -1420 359 -1380
rect 395 -1420 397 -1380
rect 511 -1380 513 -1340
rect 549 -1380 551 -1340
rect 6 -1444 46 -1442
rect 475 -1425 477 -1405
rect 1146 -1413 1148 -1373
rect 1198 -1413 1200 -1373
rect 1250 -1413 1252 -1373
rect 1302 -1413 1304 -1373
rect 1347 -1405 1349 -1365
rect 1379 -1405 1381 -1365
rect 1417 -1405 1419 -1385
rect 321 -1465 323 -1445
rect 860 -1476 862 -1436
rect 898 -1476 900 -1436
rect 1146 -1475 1148 -1435
rect 1198 -1475 1200 -1435
rect -342 -1546 -340 -1506
rect -290 -1546 -288 -1506
rect -238 -1546 -236 -1506
rect -186 -1546 -184 -1506
rect -141 -1538 -139 -1498
rect -109 -1538 -107 -1498
rect 824 -1521 826 -1501
rect -342 -1608 -340 -1568
rect -290 -1608 -288 -1568
rect 357 -1564 359 -1524
rect 395 -1564 397 -1524
rect 321 -1609 323 -1589
rect 486 -1594 488 -1554
rect 524 -1594 526 -1554
rect 450 -1639 452 -1619
rect 620 -1655 622 -1615
rect 658 -1655 660 -1615
rect 360 -1734 362 -1694
rect 398 -1734 400 -1694
rect 584 -1700 586 -1680
rect 324 -1779 326 -1759
rect 491 -1764 493 -1724
rect 529 -1764 531 -1724
rect 455 -1809 457 -1789
rect 360 -1878 362 -1838
rect 398 -1878 400 -1838
rect 749 -1844 751 -1804
rect 787 -1844 789 -1804
rect 713 -1889 715 -1869
rect 324 -1923 326 -1903
rect 360 -2005 362 -1965
rect 398 -2005 400 -1965
rect 324 -2050 326 -2030
rect 491 -2035 493 -1995
rect 529 -2035 531 -1995
rect 455 -2080 457 -2060
rect 626 -2065 628 -2025
rect 664 -2065 666 -2025
rect 360 -2149 362 -2109
rect 398 -2149 400 -2109
rect 590 -2110 592 -2090
rect 324 -2194 326 -2174
<< ndiffusion >>
rect 964 262 984 263
rect 964 259 984 260
rect 1013 252 1014 272
rect 1016 252 1017 272
rect 1013 220 1014 240
rect 1016 220 1017 240
rect 1347 264 1348 284
rect 1350 264 1351 284
rect 1379 264 1380 284
rect 1382 264 1383 284
rect 1417 274 1418 284
rect 1420 274 1421 284
rect 1250 240 1251 260
rect 1253 240 1254 260
rect 1302 240 1303 260
rect 1305 240 1306 260
rect 964 211 984 212
rect 964 208 984 209
rect 1045 193 1046 213
rect 1048 193 1049 213
rect 1146 193 1147 213
rect 1149 193 1150 213
rect 1198 193 1199 213
rect 1201 193 1202 213
rect 1250 193 1251 213
rect 1253 193 1254 213
rect 1302 193 1303 213
rect 1305 193 1306 213
rect -139 156 -138 176
rect -136 156 -135 176
rect -107 156 -106 176
rect -104 156 -103 176
rect -236 132 -235 152
rect -233 132 -232 152
rect -184 132 -183 152
rect -181 132 -180 152
rect -340 85 -339 105
rect -337 85 -336 105
rect -288 85 -287 105
rect -285 85 -284 105
rect -236 85 -235 105
rect -233 85 -232 105
rect -184 85 -183 105
rect -181 85 -180 105
rect 115 101 116 121
rect 118 101 119 121
rect 115 69 116 89
rect 118 69 119 89
rect 382 106 383 126
rect 385 106 386 126
rect 147 68 148 88
rect 150 68 151 88
rect 185 68 186 88
rect 188 68 189 88
rect 418 76 419 96
rect 421 76 422 96
rect 456 76 457 96
rect 459 76 460 96
rect 964 81 984 82
rect 964 78 984 79
rect 1013 71 1014 91
rect 1016 71 1017 91
rect 1013 39 1014 59
rect 1016 39 1017 59
rect 1346 64 1347 84
rect 1349 64 1350 84
rect 1378 64 1379 84
rect 1381 64 1382 84
rect 1416 74 1417 84
rect 1419 74 1420 84
rect 1249 40 1250 60
rect 1252 40 1253 60
rect 1301 40 1302 60
rect 1304 40 1305 60
rect 964 30 984 31
rect 66 17 86 18
rect 66 14 86 15
rect 115 7 116 27
rect 118 7 119 27
rect 115 -25 116 -5
rect 118 -25 119 -5
rect 276 -22 277 -2
rect 279 -22 280 -2
rect 964 27 984 28
rect 1045 12 1046 32
rect 1048 12 1049 32
rect 1145 -7 1146 13
rect 1148 -7 1149 13
rect 1197 -7 1198 13
rect 1200 -7 1201 13
rect 1249 -7 1250 13
rect 1252 -7 1253 13
rect 1301 -7 1302 13
rect 1304 -7 1305 13
rect 66 -34 86 -33
rect -140 -55 -139 -35
rect -137 -55 -136 -35
rect -108 -55 -107 -35
rect -105 -55 -104 -35
rect 66 -37 86 -36
rect 147 -52 148 -32
rect 150 -52 151 -32
rect 312 -52 313 -32
rect 315 -52 316 -32
rect 350 -52 351 -32
rect 353 -52 354 -32
rect -237 -79 -236 -59
rect -234 -79 -233 -59
rect -185 -79 -184 -59
rect -182 -79 -181 -59
rect -341 -126 -340 -106
rect -338 -126 -337 -106
rect -289 -126 -288 -106
rect -286 -126 -285 -106
rect -237 -126 -236 -106
rect -234 -126 -233 -106
rect -185 -126 -184 -106
rect -182 -126 -181 -106
rect 115 -189 116 -169
rect 118 -189 119 -169
rect 115 -221 116 -201
rect 118 -221 119 -201
rect 459 -184 460 -164
rect 462 -184 463 -164
rect 147 -222 148 -202
rect 150 -222 151 -202
rect 185 -222 186 -202
rect 188 -222 189 -202
rect 495 -214 496 -194
rect 498 -214 499 -194
rect 533 -214 534 -194
rect 536 -214 537 -194
rect -148 -259 -147 -239
rect -145 -259 -144 -239
rect -116 -259 -115 -239
rect -113 -259 -112 -239
rect -245 -283 -244 -263
rect -242 -283 -241 -263
rect -193 -283 -192 -263
rect -190 -283 -189 -263
rect 66 -273 86 -272
rect 66 -276 86 -275
rect 115 -283 116 -263
rect 118 -283 119 -263
rect -349 -330 -348 -310
rect -346 -330 -345 -310
rect -297 -330 -296 -310
rect -294 -330 -293 -310
rect -245 -330 -244 -310
rect -242 -330 -241 -310
rect -193 -330 -192 -310
rect -190 -330 -189 -310
rect 115 -315 116 -295
rect 118 -315 119 -295
rect 356 -312 357 -292
rect 359 -312 360 -292
rect 66 -324 86 -323
rect 66 -327 86 -326
rect 147 -342 148 -322
rect 150 -342 151 -322
rect 579 -306 580 -286
rect 582 -306 583 -286
rect 392 -342 393 -322
rect 395 -342 396 -322
rect 430 -342 431 -322
rect 433 -342 434 -322
rect 615 -336 616 -316
rect 618 -336 619 -316
rect 653 -336 654 -316
rect 656 -336 657 -316
rect 964 -331 984 -330
rect 964 -334 984 -333
rect 1013 -341 1014 -321
rect 1016 -341 1017 -321
rect 1013 -373 1014 -353
rect 1016 -373 1017 -353
rect 1345 -335 1346 -315
rect 1348 -335 1349 -315
rect 1377 -335 1378 -315
rect 1380 -335 1381 -315
rect 1415 -325 1416 -315
rect 1418 -325 1419 -315
rect 1248 -359 1249 -339
rect 1251 -359 1252 -339
rect 1300 -359 1301 -339
rect 1303 -359 1304 -339
rect 964 -382 984 -381
rect 284 -438 285 -418
rect 287 -438 288 -418
rect 964 -385 984 -384
rect 1045 -400 1046 -380
rect 1048 -400 1049 -380
rect 1144 -406 1145 -386
rect 1147 -406 1148 -386
rect 1196 -406 1197 -386
rect 1199 -406 1200 -386
rect 1248 -406 1249 -386
rect 1251 -406 1252 -386
rect 1300 -406 1301 -386
rect 1303 -406 1304 -386
rect -149 -470 -148 -450
rect -146 -470 -145 -450
rect -117 -470 -116 -450
rect -114 -470 -113 -450
rect 320 -468 321 -448
rect 323 -468 324 -448
rect 358 -468 359 -448
rect 361 -468 362 -448
rect 413 -468 414 -448
rect 416 -468 417 -448
rect -246 -494 -245 -474
rect -243 -494 -242 -474
rect -194 -494 -193 -474
rect -191 -494 -190 -474
rect 449 -498 450 -478
rect 452 -498 453 -478
rect 487 -498 488 -478
rect 490 -498 491 -478
rect -350 -541 -349 -521
rect -347 -541 -346 -521
rect -298 -541 -297 -521
rect -295 -541 -294 -521
rect -246 -541 -245 -521
rect -243 -541 -242 -521
rect -194 -541 -193 -521
rect -191 -541 -190 -521
rect 115 -606 116 -586
rect 118 -606 119 -586
rect 115 -638 116 -618
rect 118 -638 119 -618
rect 616 -601 617 -581
rect 619 -601 620 -581
rect -154 -665 -153 -645
rect -151 -665 -150 -645
rect -122 -665 -121 -645
rect -119 -665 -118 -645
rect 147 -639 148 -619
rect 150 -639 151 -619
rect 185 -639 186 -619
rect 188 -639 189 -619
rect 652 -631 653 -611
rect 655 -631 656 -611
rect 690 -631 691 -611
rect 693 -631 694 -611
rect -251 -689 -250 -669
rect -248 -689 -247 -669
rect -199 -689 -198 -669
rect -196 -689 -195 -669
rect 66 -690 86 -689
rect 66 -693 86 -692
rect 115 -700 116 -680
rect 118 -700 119 -680
rect -355 -736 -354 -716
rect -352 -736 -351 -716
rect -303 -736 -302 -716
rect -300 -736 -299 -716
rect -251 -736 -250 -716
rect -248 -736 -247 -716
rect -199 -736 -198 -716
rect -196 -736 -195 -716
rect 115 -732 116 -712
rect 118 -732 119 -712
rect 308 -729 309 -709
rect 311 -729 312 -709
rect 66 -741 86 -740
rect 66 -744 86 -743
rect 147 -759 148 -739
rect 150 -759 151 -739
rect 783 -738 784 -718
rect 786 -738 787 -718
rect 344 -759 345 -739
rect 347 -759 348 -739
rect 382 -759 383 -739
rect 385 -759 386 -739
rect 819 -768 820 -748
rect 822 -768 823 -748
rect 857 -768 858 -748
rect 860 -768 861 -748
rect 965 -763 985 -762
rect 965 -766 985 -765
rect 1014 -773 1015 -753
rect 1017 -773 1018 -753
rect 1014 -805 1015 -785
rect 1017 -805 1018 -785
rect 1345 -749 1346 -729
rect 1348 -749 1349 -729
rect 1377 -749 1378 -729
rect 1380 -749 1381 -729
rect 1415 -739 1416 -729
rect 1418 -739 1419 -729
rect 1248 -773 1249 -753
rect 1251 -773 1252 -753
rect 1300 -773 1301 -753
rect 1303 -773 1304 -753
rect 965 -814 985 -813
rect 965 -817 985 -816
rect -155 -876 -154 -856
rect -152 -876 -151 -856
rect -123 -876 -122 -856
rect -120 -876 -119 -856
rect 308 -873 309 -853
rect 311 -873 312 -853
rect 1046 -832 1047 -812
rect 1049 -832 1050 -812
rect 1144 -820 1145 -800
rect 1147 -820 1148 -800
rect 1196 -820 1197 -800
rect 1199 -820 1200 -800
rect 1248 -820 1249 -800
rect 1251 -820 1252 -800
rect 1300 -820 1301 -800
rect 1303 -820 1304 -800
rect -252 -900 -251 -880
rect -249 -900 -248 -880
rect -200 -900 -199 -880
rect -197 -900 -196 -880
rect 344 -903 345 -883
rect 347 -903 348 -883
rect 382 -903 383 -883
rect 385 -903 386 -883
rect 437 -903 438 -883
rect 440 -903 441 -883
rect -356 -947 -355 -927
rect -353 -947 -352 -927
rect -304 -947 -303 -927
rect -301 -947 -300 -927
rect -252 -947 -251 -927
rect -249 -947 -248 -927
rect -200 -947 -199 -927
rect -197 -947 -196 -927
rect 473 -933 474 -913
rect 476 -933 477 -913
rect 511 -933 512 -913
rect 514 -933 515 -913
rect 612 -957 613 -937
rect 615 -957 616 -937
rect 648 -987 649 -967
rect 651 -987 652 -967
rect 686 -987 687 -967
rect 689 -987 690 -967
rect 311 -1043 312 -1023
rect 314 -1043 315 -1023
rect 347 -1073 348 -1053
rect 350 -1073 351 -1053
rect 385 -1073 386 -1053
rect 388 -1073 389 -1053
rect 442 -1073 443 -1053
rect 445 -1073 446 -1053
rect 478 -1103 479 -1083
rect 481 -1103 482 -1083
rect 516 -1103 517 -1083
rect 519 -1103 520 -1083
rect 311 -1187 312 -1167
rect 314 -1187 315 -1167
rect 347 -1217 348 -1197
rect 350 -1217 351 -1197
rect 385 -1217 386 -1197
rect 388 -1217 389 -1197
rect 115 -1307 116 -1287
rect 118 -1307 119 -1287
rect 115 -1339 116 -1319
rect 118 -1339 119 -1319
rect -141 -1367 -140 -1347
rect -138 -1367 -137 -1347
rect -109 -1367 -108 -1347
rect -106 -1367 -105 -1347
rect 147 -1340 148 -1320
rect 150 -1340 151 -1320
rect 185 -1340 186 -1320
rect 188 -1340 189 -1320
rect -238 -1391 -237 -1371
rect -235 -1391 -234 -1371
rect -186 -1391 -185 -1371
rect -183 -1391 -182 -1371
rect 66 -1391 86 -1390
rect 66 -1394 86 -1393
rect 115 -1401 116 -1381
rect 118 -1401 119 -1381
rect -342 -1438 -341 -1418
rect -339 -1438 -338 -1418
rect -290 -1438 -289 -1418
rect -287 -1438 -286 -1418
rect -238 -1438 -237 -1418
rect -235 -1438 -234 -1418
rect -186 -1438 -185 -1418
rect -183 -1438 -182 -1418
rect 115 -1433 116 -1413
rect 118 -1433 119 -1413
rect 320 -1430 321 -1410
rect 323 -1430 324 -1410
rect 474 -1390 475 -1370
rect 477 -1390 478 -1370
rect 66 -1442 86 -1441
rect 66 -1445 86 -1444
rect 147 -1460 148 -1440
rect 150 -1460 151 -1440
rect 510 -1420 511 -1400
rect 513 -1420 514 -1400
rect 548 -1420 549 -1400
rect 551 -1420 552 -1400
rect 356 -1460 357 -1440
rect 359 -1460 360 -1440
rect 394 -1460 395 -1440
rect 397 -1460 398 -1440
rect 823 -1486 824 -1466
rect 826 -1486 827 -1466
rect 1346 -1445 1347 -1425
rect 1349 -1445 1350 -1425
rect 1378 -1445 1379 -1425
rect 1381 -1445 1382 -1425
rect 1416 -1435 1417 -1425
rect 1419 -1435 1420 -1425
rect 1249 -1469 1250 -1449
rect 1252 -1469 1253 -1449
rect 1301 -1469 1302 -1449
rect 1304 -1469 1305 -1449
rect 859 -1516 860 -1496
rect 862 -1516 863 -1496
rect 897 -1516 898 -1496
rect 900 -1516 901 -1496
rect 1145 -1516 1146 -1496
rect 1148 -1516 1149 -1496
rect 1197 -1516 1198 -1496
rect 1200 -1516 1201 -1496
rect 1249 -1516 1250 -1496
rect 1252 -1516 1253 -1496
rect 1301 -1516 1302 -1496
rect 1304 -1516 1305 -1496
rect -142 -1578 -141 -1558
rect -139 -1578 -138 -1558
rect -110 -1578 -109 -1558
rect -107 -1578 -106 -1558
rect 320 -1574 321 -1554
rect 323 -1574 324 -1554
rect -239 -1602 -238 -1582
rect -236 -1602 -235 -1582
rect -187 -1602 -186 -1582
rect -184 -1602 -183 -1582
rect 356 -1604 357 -1584
rect 359 -1604 360 -1584
rect 394 -1604 395 -1584
rect 397 -1604 398 -1584
rect 449 -1604 450 -1584
rect 452 -1604 453 -1584
rect -343 -1649 -342 -1629
rect -340 -1649 -339 -1629
rect -291 -1649 -290 -1629
rect -288 -1649 -287 -1629
rect -239 -1649 -238 -1629
rect -236 -1649 -235 -1629
rect -187 -1649 -186 -1629
rect -184 -1649 -183 -1629
rect 485 -1634 486 -1614
rect 488 -1634 489 -1614
rect 523 -1634 524 -1614
rect 526 -1634 527 -1614
rect 583 -1665 584 -1645
rect 586 -1665 587 -1645
rect 323 -1744 324 -1724
rect 326 -1744 327 -1724
rect 619 -1695 620 -1675
rect 622 -1695 623 -1675
rect 657 -1695 658 -1675
rect 660 -1695 661 -1675
rect 359 -1774 360 -1754
rect 362 -1774 363 -1754
rect 397 -1774 398 -1754
rect 400 -1774 401 -1754
rect 454 -1774 455 -1754
rect 457 -1774 458 -1754
rect 490 -1804 491 -1784
rect 493 -1804 494 -1784
rect 528 -1804 529 -1784
rect 531 -1804 532 -1784
rect 323 -1888 324 -1868
rect 326 -1888 327 -1868
rect 712 -1854 713 -1834
rect 715 -1854 716 -1834
rect 748 -1884 749 -1864
rect 751 -1884 752 -1864
rect 786 -1884 787 -1864
rect 789 -1884 790 -1864
rect 359 -1918 360 -1898
rect 362 -1918 363 -1898
rect 397 -1918 398 -1898
rect 400 -1918 401 -1898
rect 323 -2015 324 -1995
rect 326 -2015 327 -1995
rect 359 -2045 360 -2025
rect 362 -2045 363 -2025
rect 397 -2045 398 -2025
rect 400 -2045 401 -2025
rect 454 -2045 455 -2025
rect 457 -2045 458 -2025
rect 490 -2075 491 -2055
rect 493 -2075 494 -2055
rect 528 -2075 529 -2055
rect 531 -2075 532 -2055
rect 589 -2075 590 -2055
rect 592 -2075 593 -2055
rect 323 -2159 324 -2139
rect 326 -2159 327 -2139
rect 625 -2105 626 -2085
rect 628 -2105 629 -2085
rect 663 -2105 664 -2085
rect 666 -2105 667 -2085
rect 359 -2189 360 -2169
rect 362 -2189 363 -2169
rect 397 -2189 398 -2169
rect 400 -2189 401 -2169
<< pdiffusion >>
rect 1146 296 1147 336
rect 1149 296 1150 336
rect 1198 296 1199 336
rect 1201 296 1202 336
rect 1250 296 1251 336
rect 1253 296 1254 336
rect 1302 296 1303 336
rect 1305 296 1306 336
rect 1347 304 1348 344
rect 1350 304 1351 344
rect 1379 304 1380 344
rect 1382 304 1383 344
rect 1417 304 1418 324
rect 1420 304 1421 324
rect 904 262 944 263
rect 904 259 944 260
rect -340 188 -339 228
rect -337 188 -336 228
rect -288 188 -287 228
rect -285 188 -284 228
rect -236 188 -235 228
rect -233 188 -232 228
rect -184 188 -183 228
rect -181 188 -180 228
rect -139 196 -138 236
rect -136 196 -135 236
rect -107 196 -106 236
rect -104 196 -103 236
rect 1045 233 1046 273
rect 1048 233 1049 273
rect 1146 234 1147 274
rect 1149 234 1150 274
rect 1198 234 1199 274
rect 1201 234 1202 274
rect 904 211 944 212
rect 904 208 944 209
rect -340 126 -339 166
rect -337 126 -336 166
rect -288 126 -287 166
rect -285 126 -284 166
rect 147 108 148 148
rect 150 108 151 148
rect 185 108 186 148
rect 188 108 189 148
rect 418 116 419 156
rect 421 116 422 156
rect 456 116 457 156
rect 459 116 460 156
rect 382 71 383 91
rect 385 71 386 91
rect 1145 96 1146 136
rect 1148 96 1149 136
rect 1197 96 1198 136
rect 1200 96 1201 136
rect 1249 96 1250 136
rect 1252 96 1253 136
rect 1301 96 1302 136
rect 1304 96 1305 136
rect 1346 104 1347 144
rect 1349 104 1350 144
rect 1378 104 1379 144
rect 1381 104 1382 144
rect 1416 104 1417 124
rect 1419 104 1420 124
rect 904 81 944 82
rect 904 78 944 79
rect 1045 52 1046 92
rect 1048 52 1049 92
rect 904 30 944 31
rect 1145 34 1146 74
rect 1148 34 1149 74
rect 1197 34 1198 74
rect 1200 34 1201 74
rect -341 -23 -340 17
rect -338 -23 -337 17
rect -289 -23 -288 17
rect -286 -23 -285 17
rect -237 -23 -236 17
rect -234 -23 -233 17
rect -185 -23 -184 17
rect -182 -23 -181 17
rect -140 -15 -139 25
rect -137 -15 -136 25
rect -108 -15 -107 25
rect -105 -15 -104 25
rect 6 17 46 18
rect 6 14 46 15
rect 147 -12 148 28
rect 150 -12 151 28
rect 6 -34 46 -33
rect 312 -12 313 28
rect 315 -12 316 28
rect 350 -12 351 28
rect 353 -12 354 28
rect 904 27 944 28
rect -341 -85 -340 -45
rect -338 -85 -337 -45
rect -289 -85 -288 -45
rect -286 -85 -285 -45
rect 6 -37 46 -36
rect 276 -57 277 -37
rect 279 -57 280 -37
rect -349 -227 -348 -187
rect -346 -227 -345 -187
rect -297 -227 -296 -187
rect -294 -227 -293 -187
rect -245 -227 -244 -187
rect -242 -227 -241 -187
rect -193 -227 -192 -187
rect -190 -227 -189 -187
rect -148 -219 -147 -179
rect -145 -219 -144 -179
rect -116 -219 -115 -179
rect -113 -219 -112 -179
rect 147 -182 148 -142
rect 150 -182 151 -142
rect 185 -182 186 -142
rect 188 -182 189 -142
rect 495 -174 496 -134
rect 498 -174 499 -134
rect 533 -174 534 -134
rect 536 -174 537 -134
rect 459 -219 460 -199
rect 462 -219 463 -199
rect -349 -289 -348 -249
rect -346 -289 -345 -249
rect -297 -289 -296 -249
rect -294 -289 -293 -249
rect 6 -273 46 -272
rect 6 -276 46 -275
rect 147 -302 148 -262
rect 150 -302 151 -262
rect 6 -324 46 -323
rect 392 -302 393 -262
rect 395 -302 396 -262
rect 430 -302 431 -262
rect 433 -302 434 -262
rect 6 -327 46 -326
rect 615 -296 616 -256
rect 618 -296 619 -256
rect 653 -296 654 -256
rect 656 -296 657 -256
rect 1144 -303 1145 -263
rect 1147 -303 1148 -263
rect 1196 -303 1197 -263
rect 1199 -303 1200 -263
rect 1248 -303 1249 -263
rect 1251 -303 1252 -263
rect 1300 -303 1301 -263
rect 1303 -303 1304 -263
rect 1345 -295 1346 -255
rect 1348 -295 1349 -255
rect 1377 -295 1378 -255
rect 1380 -295 1381 -255
rect 1415 -295 1416 -275
rect 1418 -295 1419 -275
rect 356 -347 357 -327
rect 359 -347 360 -327
rect 579 -341 580 -321
rect 582 -341 583 -321
rect 904 -331 944 -330
rect 904 -334 944 -333
rect 1045 -360 1046 -320
rect 1048 -360 1049 -320
rect 904 -382 944 -381
rect 1144 -365 1145 -325
rect 1147 -365 1148 -325
rect 1196 -365 1197 -325
rect 1199 -365 1200 -325
rect 904 -385 944 -384
rect -350 -438 -349 -398
rect -347 -438 -346 -398
rect -298 -438 -297 -398
rect -295 -438 -294 -398
rect -246 -438 -245 -398
rect -243 -438 -242 -398
rect -194 -438 -193 -398
rect -191 -438 -190 -398
rect -149 -430 -148 -390
rect -146 -430 -145 -390
rect -117 -430 -116 -390
rect -114 -430 -113 -390
rect 320 -428 321 -388
rect 323 -428 324 -388
rect 358 -428 359 -388
rect 361 -428 362 -388
rect -350 -500 -349 -460
rect -347 -500 -346 -460
rect -298 -500 -297 -460
rect -295 -500 -294 -460
rect 284 -473 285 -453
rect 287 -473 288 -453
rect 449 -458 450 -418
rect 452 -458 453 -418
rect 487 -458 488 -418
rect 490 -458 491 -418
rect 413 -503 414 -483
rect 416 -503 417 -483
rect -355 -633 -354 -593
rect -352 -633 -351 -593
rect -303 -633 -302 -593
rect -300 -633 -299 -593
rect -251 -633 -250 -593
rect -248 -633 -247 -593
rect -199 -633 -198 -593
rect -196 -633 -195 -593
rect -154 -625 -153 -585
rect -151 -625 -150 -585
rect -122 -625 -121 -585
rect -119 -625 -118 -585
rect 147 -599 148 -559
rect 150 -599 151 -559
rect 185 -599 186 -559
rect 188 -599 189 -559
rect 652 -591 653 -551
rect 655 -591 656 -551
rect 690 -591 691 -551
rect 693 -591 694 -551
rect -355 -695 -354 -655
rect -352 -695 -351 -655
rect -303 -695 -302 -655
rect -300 -695 -299 -655
rect 616 -636 617 -616
rect 619 -636 620 -616
rect 6 -690 46 -689
rect 6 -693 46 -692
rect 147 -719 148 -679
rect 150 -719 151 -679
rect 6 -741 46 -740
rect 344 -719 345 -679
rect 347 -719 348 -679
rect 382 -719 383 -679
rect 385 -719 386 -679
rect 6 -744 46 -743
rect 819 -728 820 -688
rect 822 -728 823 -688
rect 857 -728 858 -688
rect 860 -728 861 -688
rect 1144 -717 1145 -677
rect 1147 -717 1148 -677
rect 1196 -717 1197 -677
rect 1199 -717 1200 -677
rect 1248 -717 1249 -677
rect 1251 -717 1252 -677
rect 1300 -717 1301 -677
rect 1303 -717 1304 -677
rect 1345 -709 1346 -669
rect 1348 -709 1349 -669
rect 1377 -709 1378 -669
rect 1380 -709 1381 -669
rect 1415 -709 1416 -689
rect 1418 -709 1419 -689
rect 308 -764 309 -744
rect 311 -764 312 -744
rect 783 -773 784 -753
rect 786 -773 787 -753
rect 905 -763 945 -762
rect 905 -766 945 -765
rect -356 -844 -355 -804
rect -353 -844 -352 -804
rect -304 -844 -303 -804
rect -301 -844 -300 -804
rect -252 -844 -251 -804
rect -249 -844 -248 -804
rect -200 -844 -199 -804
rect -197 -844 -196 -804
rect -155 -836 -154 -796
rect -152 -836 -151 -796
rect -123 -836 -122 -796
rect -120 -836 -119 -796
rect 1046 -792 1047 -752
rect 1049 -792 1050 -752
rect 1144 -779 1145 -739
rect 1147 -779 1148 -739
rect 1196 -779 1197 -739
rect 1199 -779 1200 -739
rect 905 -814 945 -813
rect 905 -817 945 -816
rect -356 -906 -355 -866
rect -353 -906 -352 -866
rect -304 -906 -303 -866
rect -301 -906 -300 -866
rect 344 -863 345 -823
rect 347 -863 348 -823
rect 382 -863 383 -823
rect 385 -863 386 -823
rect 308 -908 309 -888
rect 311 -908 312 -888
rect 473 -893 474 -853
rect 476 -893 477 -853
rect 511 -893 512 -853
rect 514 -893 515 -853
rect 437 -938 438 -918
rect 440 -938 441 -918
rect 648 -947 649 -907
rect 651 -947 652 -907
rect 686 -947 687 -907
rect 689 -947 690 -907
rect 612 -992 613 -972
rect 615 -992 616 -972
rect 347 -1033 348 -993
rect 350 -1033 351 -993
rect 385 -1033 386 -993
rect 388 -1033 389 -993
rect 311 -1078 312 -1058
rect 314 -1078 315 -1058
rect 478 -1063 479 -1023
rect 481 -1063 482 -1023
rect 516 -1063 517 -1023
rect 519 -1063 520 -1023
rect 442 -1108 443 -1088
rect 445 -1108 446 -1088
rect 347 -1177 348 -1137
rect 350 -1177 351 -1137
rect 385 -1177 386 -1137
rect 388 -1177 389 -1137
rect 311 -1222 312 -1202
rect 314 -1222 315 -1202
rect -342 -1335 -341 -1295
rect -339 -1335 -338 -1295
rect -290 -1335 -289 -1295
rect -287 -1335 -286 -1295
rect -238 -1335 -237 -1295
rect -235 -1335 -234 -1295
rect -186 -1335 -185 -1295
rect -183 -1335 -182 -1295
rect -141 -1327 -140 -1287
rect -138 -1327 -137 -1287
rect -109 -1327 -108 -1287
rect -106 -1327 -105 -1287
rect 147 -1300 148 -1260
rect 150 -1300 151 -1260
rect 185 -1300 186 -1260
rect 188 -1300 189 -1260
rect -342 -1397 -341 -1357
rect -339 -1397 -338 -1357
rect -290 -1397 -289 -1357
rect -287 -1397 -286 -1357
rect 6 -1391 46 -1390
rect 6 -1394 46 -1393
rect 147 -1420 148 -1380
rect 150 -1420 151 -1380
rect 6 -1442 46 -1441
rect 356 -1420 357 -1380
rect 359 -1420 360 -1380
rect 394 -1420 395 -1380
rect 397 -1420 398 -1380
rect 510 -1380 511 -1340
rect 513 -1380 514 -1340
rect 548 -1380 549 -1340
rect 551 -1380 552 -1340
rect 6 -1445 46 -1444
rect 474 -1425 475 -1405
rect 477 -1425 478 -1405
rect 1145 -1413 1146 -1373
rect 1148 -1413 1149 -1373
rect 1197 -1413 1198 -1373
rect 1200 -1413 1201 -1373
rect 1249 -1413 1250 -1373
rect 1252 -1413 1253 -1373
rect 1301 -1413 1302 -1373
rect 1304 -1413 1305 -1373
rect 1346 -1405 1347 -1365
rect 1349 -1405 1350 -1365
rect 1378 -1405 1379 -1365
rect 1381 -1405 1382 -1365
rect 1416 -1405 1417 -1385
rect 1419 -1405 1420 -1385
rect 320 -1465 321 -1445
rect 323 -1465 324 -1445
rect 859 -1476 860 -1436
rect 862 -1476 863 -1436
rect 897 -1476 898 -1436
rect 900 -1476 901 -1436
rect 1145 -1475 1146 -1435
rect 1148 -1475 1149 -1435
rect 1197 -1475 1198 -1435
rect 1200 -1475 1201 -1435
rect -343 -1546 -342 -1506
rect -340 -1546 -339 -1506
rect -291 -1546 -290 -1506
rect -288 -1546 -287 -1506
rect -239 -1546 -238 -1506
rect -236 -1546 -235 -1506
rect -187 -1546 -186 -1506
rect -184 -1546 -183 -1506
rect -142 -1538 -141 -1498
rect -139 -1538 -138 -1498
rect -110 -1538 -109 -1498
rect -107 -1538 -106 -1498
rect 823 -1521 824 -1501
rect 826 -1521 827 -1501
rect -343 -1608 -342 -1568
rect -340 -1608 -339 -1568
rect -291 -1608 -290 -1568
rect -288 -1608 -287 -1568
rect 356 -1564 357 -1524
rect 359 -1564 360 -1524
rect 394 -1564 395 -1524
rect 397 -1564 398 -1524
rect 320 -1609 321 -1589
rect 323 -1609 324 -1589
rect 485 -1594 486 -1554
rect 488 -1594 489 -1554
rect 523 -1594 524 -1554
rect 526 -1594 527 -1554
rect 449 -1639 450 -1619
rect 452 -1639 453 -1619
rect 619 -1655 620 -1615
rect 622 -1655 623 -1615
rect 657 -1655 658 -1615
rect 660 -1655 661 -1615
rect 359 -1734 360 -1694
rect 362 -1734 363 -1694
rect 397 -1734 398 -1694
rect 400 -1734 401 -1694
rect 583 -1700 584 -1680
rect 586 -1700 587 -1680
rect 323 -1779 324 -1759
rect 326 -1779 327 -1759
rect 490 -1764 491 -1724
rect 493 -1764 494 -1724
rect 528 -1764 529 -1724
rect 531 -1764 532 -1724
rect 454 -1809 455 -1789
rect 457 -1809 458 -1789
rect 359 -1878 360 -1838
rect 362 -1878 363 -1838
rect 397 -1878 398 -1838
rect 400 -1878 401 -1838
rect 748 -1844 749 -1804
rect 751 -1844 752 -1804
rect 786 -1844 787 -1804
rect 789 -1844 790 -1804
rect 712 -1889 713 -1869
rect 715 -1889 716 -1869
rect 323 -1923 324 -1903
rect 326 -1923 327 -1903
rect 359 -2005 360 -1965
rect 362 -2005 363 -1965
rect 397 -2005 398 -1965
rect 400 -2005 401 -1965
rect 323 -2050 324 -2030
rect 326 -2050 327 -2030
rect 490 -2035 491 -1995
rect 493 -2035 494 -1995
rect 528 -2035 529 -1995
rect 531 -2035 532 -1995
rect 454 -2080 455 -2060
rect 457 -2080 458 -2060
rect 625 -2065 626 -2025
rect 628 -2065 629 -2025
rect 663 -2065 664 -2025
rect 666 -2065 667 -2025
rect 359 -2149 360 -2109
rect 362 -2149 363 -2109
rect 397 -2149 398 -2109
rect 400 -2149 401 -2109
rect 589 -2110 590 -2090
rect 592 -2110 593 -2090
rect 323 -2194 324 -2174
rect 326 -2194 327 -2174
<< ndcontact >>
rect 964 263 984 267
rect 964 255 984 259
rect 1009 252 1013 272
rect 1017 252 1021 272
rect 1009 220 1013 240
rect 1017 220 1021 240
rect 1343 264 1347 284
rect 1351 264 1355 284
rect 1375 264 1379 284
rect 1383 264 1387 284
rect 1413 274 1417 284
rect 1421 274 1425 284
rect 1246 240 1250 260
rect 1254 240 1258 260
rect 1298 240 1302 260
rect 1306 240 1310 260
rect 964 212 984 216
rect 964 204 984 208
rect 1041 193 1045 213
rect 1049 193 1053 213
rect 1142 193 1146 213
rect 1150 193 1154 213
rect 1194 193 1198 213
rect 1202 193 1206 213
rect 1246 193 1250 213
rect 1254 193 1258 213
rect 1298 193 1302 213
rect 1306 193 1310 213
rect -143 156 -139 176
rect -135 156 -131 176
rect -111 156 -107 176
rect -103 156 -99 176
rect -240 132 -236 152
rect -232 132 -228 152
rect -188 132 -184 152
rect -180 132 -176 152
rect -344 85 -340 105
rect -336 85 -332 105
rect -292 85 -288 105
rect -284 85 -280 105
rect -240 85 -236 105
rect -232 85 -228 105
rect -188 85 -184 105
rect -180 85 -176 105
rect 111 101 115 121
rect 119 101 123 121
rect 111 69 115 89
rect 119 69 123 89
rect 378 106 382 126
rect 386 106 390 126
rect 143 68 147 88
rect 151 68 155 88
rect 181 68 185 88
rect 189 68 193 88
rect 414 76 418 96
rect 422 76 426 96
rect 452 76 456 96
rect 460 76 464 96
rect 964 82 984 86
rect 964 74 984 78
rect 1009 71 1013 91
rect 1017 71 1021 91
rect 1009 39 1013 59
rect 1017 39 1021 59
rect 964 31 984 35
rect 1342 64 1346 84
rect 1350 64 1354 84
rect 1374 64 1378 84
rect 1382 64 1386 84
rect 1412 74 1416 84
rect 1420 74 1424 84
rect 1245 40 1249 60
rect 1253 40 1257 60
rect 1297 40 1301 60
rect 1305 40 1309 60
rect 66 18 86 22
rect 66 10 86 14
rect 111 7 115 27
rect 119 7 123 27
rect 111 -25 115 -5
rect 119 -25 123 -5
rect 66 -33 86 -29
rect 272 -22 276 -2
rect 280 -22 284 -2
rect 964 23 984 27
rect 1041 12 1045 32
rect 1049 12 1053 32
rect 1141 -7 1145 13
rect 1149 -7 1153 13
rect 1193 -7 1197 13
rect 1201 -7 1205 13
rect 1245 -7 1249 13
rect 1253 -7 1257 13
rect 1297 -7 1301 13
rect 1305 -7 1309 13
rect -144 -55 -140 -35
rect -136 -55 -132 -35
rect -112 -55 -108 -35
rect -104 -55 -100 -35
rect 66 -41 86 -37
rect 143 -52 147 -32
rect 151 -52 155 -32
rect 308 -52 312 -32
rect 316 -52 320 -32
rect 346 -52 350 -32
rect 354 -52 358 -32
rect -241 -79 -237 -59
rect -233 -79 -229 -59
rect -189 -79 -185 -59
rect -181 -79 -177 -59
rect -345 -126 -341 -106
rect -337 -126 -333 -106
rect -293 -126 -289 -106
rect -285 -126 -281 -106
rect -241 -126 -237 -106
rect -233 -126 -229 -106
rect -189 -126 -185 -106
rect -181 -126 -177 -106
rect 111 -189 115 -169
rect 119 -189 123 -169
rect 111 -221 115 -201
rect 119 -221 123 -201
rect 455 -184 459 -164
rect 463 -184 467 -164
rect 143 -222 147 -202
rect 151 -222 155 -202
rect 181 -222 185 -202
rect 189 -222 193 -202
rect 491 -214 495 -194
rect 499 -214 503 -194
rect 529 -214 533 -194
rect 537 -214 541 -194
rect -152 -259 -148 -239
rect -144 -259 -140 -239
rect -120 -259 -116 -239
rect -112 -259 -108 -239
rect -249 -283 -245 -263
rect -241 -283 -237 -263
rect -197 -283 -193 -263
rect -189 -283 -185 -263
rect 66 -272 86 -268
rect 66 -280 86 -276
rect 111 -283 115 -263
rect 119 -283 123 -263
rect -353 -330 -349 -310
rect -345 -330 -341 -310
rect -301 -330 -297 -310
rect -293 -330 -289 -310
rect -249 -330 -245 -310
rect -241 -330 -237 -310
rect -197 -330 -193 -310
rect -189 -330 -185 -310
rect 111 -315 115 -295
rect 119 -315 123 -295
rect 66 -323 86 -319
rect 352 -312 356 -292
rect 360 -312 364 -292
rect 66 -331 86 -327
rect 143 -342 147 -322
rect 151 -342 155 -322
rect 575 -306 579 -286
rect 583 -306 587 -286
rect 388 -342 392 -322
rect 396 -342 400 -322
rect 426 -342 430 -322
rect 434 -342 438 -322
rect 611 -336 615 -316
rect 619 -336 623 -316
rect 649 -336 653 -316
rect 657 -336 661 -316
rect 964 -330 984 -326
rect 964 -338 984 -334
rect 1009 -341 1013 -321
rect 1017 -341 1021 -321
rect 1009 -373 1013 -353
rect 1017 -373 1021 -353
rect 964 -381 984 -377
rect 1341 -335 1345 -315
rect 1349 -335 1353 -315
rect 1373 -335 1377 -315
rect 1381 -335 1385 -315
rect 1411 -325 1415 -315
rect 1419 -325 1423 -315
rect 1244 -359 1248 -339
rect 1252 -359 1256 -339
rect 1296 -359 1300 -339
rect 1304 -359 1308 -339
rect 280 -438 284 -418
rect 288 -438 292 -418
rect 964 -389 984 -385
rect 1041 -400 1045 -380
rect 1049 -400 1053 -380
rect 1140 -406 1144 -386
rect 1148 -406 1152 -386
rect 1192 -406 1196 -386
rect 1200 -406 1204 -386
rect 1244 -406 1248 -386
rect 1252 -406 1256 -386
rect 1296 -406 1300 -386
rect 1304 -406 1308 -386
rect -153 -470 -149 -450
rect -145 -470 -141 -450
rect -121 -470 -117 -450
rect -113 -470 -109 -450
rect 316 -468 320 -448
rect 324 -468 328 -448
rect 354 -468 358 -448
rect 362 -468 366 -448
rect 409 -468 413 -448
rect 417 -468 421 -448
rect -250 -494 -246 -474
rect -242 -494 -238 -474
rect -198 -494 -194 -474
rect -190 -494 -186 -474
rect 445 -498 449 -478
rect 453 -498 457 -478
rect 483 -498 487 -478
rect 491 -498 495 -478
rect -354 -541 -350 -521
rect -346 -541 -342 -521
rect -302 -541 -298 -521
rect -294 -541 -290 -521
rect -250 -541 -246 -521
rect -242 -541 -238 -521
rect -198 -541 -194 -521
rect -190 -541 -186 -521
rect 111 -606 115 -586
rect 119 -606 123 -586
rect 111 -638 115 -618
rect 119 -638 123 -618
rect 612 -601 616 -581
rect 620 -601 624 -581
rect -158 -665 -154 -645
rect -150 -665 -146 -645
rect -126 -665 -122 -645
rect -118 -665 -114 -645
rect 143 -639 147 -619
rect 151 -639 155 -619
rect 181 -639 185 -619
rect 189 -639 193 -619
rect 648 -631 652 -611
rect 656 -631 660 -611
rect 686 -631 690 -611
rect 694 -631 698 -611
rect -255 -689 -251 -669
rect -247 -689 -243 -669
rect -203 -689 -199 -669
rect -195 -689 -191 -669
rect 66 -689 86 -685
rect 66 -697 86 -693
rect 111 -700 115 -680
rect 119 -700 123 -680
rect -359 -736 -355 -716
rect -351 -736 -347 -716
rect -307 -736 -303 -716
rect -299 -736 -295 -716
rect -255 -736 -251 -716
rect -247 -736 -243 -716
rect -203 -736 -199 -716
rect -195 -736 -191 -716
rect 111 -732 115 -712
rect 119 -732 123 -712
rect 66 -740 86 -736
rect 304 -729 308 -709
rect 312 -729 316 -709
rect 66 -748 86 -744
rect 143 -759 147 -739
rect 151 -759 155 -739
rect 779 -738 783 -718
rect 787 -738 791 -718
rect 340 -759 344 -739
rect 348 -759 352 -739
rect 378 -759 382 -739
rect 386 -759 390 -739
rect 815 -768 819 -748
rect 823 -768 827 -748
rect 853 -768 857 -748
rect 861 -768 865 -748
rect 965 -762 985 -758
rect 965 -770 985 -766
rect 1010 -773 1014 -753
rect 1018 -773 1022 -753
rect 1010 -805 1014 -785
rect 1018 -805 1022 -785
rect 1341 -749 1345 -729
rect 1349 -749 1353 -729
rect 1373 -749 1377 -729
rect 1381 -749 1385 -729
rect 1411 -739 1415 -729
rect 1419 -739 1423 -729
rect 1244 -773 1248 -753
rect 1252 -773 1256 -753
rect 1296 -773 1300 -753
rect 1304 -773 1308 -753
rect 965 -813 985 -809
rect 965 -821 985 -817
rect -159 -876 -155 -856
rect -151 -876 -147 -856
rect -127 -876 -123 -856
rect -119 -876 -115 -856
rect 304 -873 308 -853
rect 312 -873 316 -853
rect 1042 -832 1046 -812
rect 1050 -832 1054 -812
rect 1140 -820 1144 -800
rect 1148 -820 1152 -800
rect 1192 -820 1196 -800
rect 1200 -820 1204 -800
rect 1244 -820 1248 -800
rect 1252 -820 1256 -800
rect 1296 -820 1300 -800
rect 1304 -820 1308 -800
rect -256 -900 -252 -880
rect -248 -900 -244 -880
rect -204 -900 -200 -880
rect -196 -900 -192 -880
rect 340 -903 344 -883
rect 348 -903 352 -883
rect 378 -903 382 -883
rect 386 -903 390 -883
rect 433 -903 437 -883
rect 441 -903 445 -883
rect -360 -947 -356 -927
rect -352 -947 -348 -927
rect -308 -947 -304 -927
rect -300 -947 -296 -927
rect -256 -947 -252 -927
rect -248 -947 -244 -927
rect -204 -947 -200 -927
rect -196 -947 -192 -927
rect 469 -933 473 -913
rect 477 -933 481 -913
rect 507 -933 511 -913
rect 515 -933 519 -913
rect 608 -957 612 -937
rect 616 -957 620 -937
rect 644 -987 648 -967
rect 652 -987 656 -967
rect 682 -987 686 -967
rect 690 -987 694 -967
rect 307 -1043 311 -1023
rect 315 -1043 319 -1023
rect 343 -1073 347 -1053
rect 351 -1073 355 -1053
rect 381 -1073 385 -1053
rect 389 -1073 393 -1053
rect 438 -1073 442 -1053
rect 446 -1073 450 -1053
rect 474 -1103 478 -1083
rect 482 -1103 486 -1083
rect 512 -1103 516 -1083
rect 520 -1103 524 -1083
rect 307 -1187 311 -1167
rect 315 -1187 319 -1167
rect 343 -1217 347 -1197
rect 351 -1217 355 -1197
rect 381 -1217 385 -1197
rect 389 -1217 393 -1197
rect 111 -1307 115 -1287
rect 119 -1307 123 -1287
rect 111 -1339 115 -1319
rect 119 -1339 123 -1319
rect -145 -1367 -141 -1347
rect -137 -1367 -133 -1347
rect -113 -1367 -109 -1347
rect -105 -1367 -101 -1347
rect 143 -1340 147 -1320
rect 151 -1340 155 -1320
rect 181 -1340 185 -1320
rect 189 -1340 193 -1320
rect -242 -1391 -238 -1371
rect -234 -1391 -230 -1371
rect -190 -1391 -186 -1371
rect -182 -1391 -178 -1371
rect 66 -1390 86 -1386
rect 66 -1398 86 -1394
rect 111 -1401 115 -1381
rect 119 -1401 123 -1381
rect -346 -1438 -342 -1418
rect -338 -1438 -334 -1418
rect -294 -1438 -290 -1418
rect -286 -1438 -282 -1418
rect -242 -1438 -238 -1418
rect -234 -1438 -230 -1418
rect -190 -1438 -186 -1418
rect -182 -1438 -178 -1418
rect 111 -1433 115 -1413
rect 119 -1433 123 -1413
rect 66 -1441 86 -1437
rect 316 -1430 320 -1410
rect 324 -1430 328 -1410
rect 470 -1390 474 -1370
rect 478 -1390 482 -1370
rect 66 -1449 86 -1445
rect 143 -1460 147 -1440
rect 151 -1460 155 -1440
rect 506 -1420 510 -1400
rect 514 -1420 518 -1400
rect 544 -1420 548 -1400
rect 552 -1420 556 -1400
rect 352 -1460 356 -1440
rect 360 -1460 364 -1440
rect 390 -1460 394 -1440
rect 398 -1460 402 -1440
rect 819 -1486 823 -1466
rect 827 -1486 831 -1466
rect 1342 -1445 1346 -1425
rect 1350 -1445 1354 -1425
rect 1374 -1445 1378 -1425
rect 1382 -1445 1386 -1425
rect 1412 -1435 1416 -1425
rect 1420 -1435 1424 -1425
rect 1245 -1469 1249 -1449
rect 1253 -1469 1257 -1449
rect 1297 -1469 1301 -1449
rect 1305 -1469 1309 -1449
rect 855 -1516 859 -1496
rect 863 -1516 867 -1496
rect 893 -1516 897 -1496
rect 901 -1516 905 -1496
rect 1141 -1516 1145 -1496
rect 1149 -1516 1153 -1496
rect 1193 -1516 1197 -1496
rect 1201 -1516 1205 -1496
rect 1245 -1516 1249 -1496
rect 1253 -1516 1257 -1496
rect 1297 -1516 1301 -1496
rect 1305 -1516 1309 -1496
rect -146 -1578 -142 -1558
rect -138 -1578 -134 -1558
rect -114 -1578 -110 -1558
rect -106 -1578 -102 -1558
rect 316 -1574 320 -1554
rect 324 -1574 328 -1554
rect -243 -1602 -239 -1582
rect -235 -1602 -231 -1582
rect -191 -1602 -187 -1582
rect -183 -1602 -179 -1582
rect 352 -1604 356 -1584
rect 360 -1604 364 -1584
rect 390 -1604 394 -1584
rect 398 -1604 402 -1584
rect 445 -1604 449 -1584
rect 453 -1604 457 -1584
rect -347 -1649 -343 -1629
rect -339 -1649 -335 -1629
rect -295 -1649 -291 -1629
rect -287 -1649 -283 -1629
rect -243 -1649 -239 -1629
rect -235 -1649 -231 -1629
rect -191 -1649 -187 -1629
rect -183 -1649 -179 -1629
rect 481 -1634 485 -1614
rect 489 -1634 493 -1614
rect 519 -1634 523 -1614
rect 527 -1634 531 -1614
rect 579 -1665 583 -1645
rect 587 -1665 591 -1645
rect 319 -1744 323 -1724
rect 327 -1744 331 -1724
rect 615 -1695 619 -1675
rect 623 -1695 627 -1675
rect 653 -1695 657 -1675
rect 661 -1695 665 -1675
rect 355 -1774 359 -1754
rect 363 -1774 367 -1754
rect 393 -1774 397 -1754
rect 401 -1774 405 -1754
rect 450 -1774 454 -1754
rect 458 -1774 462 -1754
rect 486 -1804 490 -1784
rect 494 -1804 498 -1784
rect 524 -1804 528 -1784
rect 532 -1804 536 -1784
rect 319 -1888 323 -1868
rect 327 -1888 331 -1868
rect 708 -1854 712 -1834
rect 716 -1854 720 -1834
rect 744 -1884 748 -1864
rect 752 -1884 756 -1864
rect 782 -1884 786 -1864
rect 790 -1884 794 -1864
rect 355 -1918 359 -1898
rect 363 -1918 367 -1898
rect 393 -1918 397 -1898
rect 401 -1918 405 -1898
rect 319 -2015 323 -1995
rect 327 -2015 331 -1995
rect 355 -2045 359 -2025
rect 363 -2045 367 -2025
rect 393 -2045 397 -2025
rect 401 -2045 405 -2025
rect 450 -2045 454 -2025
rect 458 -2045 462 -2025
rect 486 -2075 490 -2055
rect 494 -2075 498 -2055
rect 524 -2075 528 -2055
rect 532 -2075 536 -2055
rect 585 -2075 589 -2055
rect 593 -2075 597 -2055
rect 319 -2159 323 -2139
rect 327 -2159 331 -2139
rect 621 -2105 625 -2085
rect 629 -2105 633 -2085
rect 659 -2105 663 -2085
rect 667 -2105 671 -2085
rect 355 -2189 359 -2169
rect 363 -2189 367 -2169
rect 393 -2189 397 -2169
rect 401 -2189 405 -2169
<< pdcontact >>
rect 1142 296 1146 336
rect 1150 296 1154 336
rect 1194 296 1198 336
rect 1202 296 1206 336
rect 1246 296 1250 336
rect 1254 296 1258 336
rect 1298 296 1302 336
rect 1306 296 1310 336
rect 1343 304 1347 344
rect 1351 304 1355 344
rect 1375 304 1379 344
rect 1383 304 1387 344
rect 1413 304 1417 324
rect 1421 304 1425 324
rect 904 263 944 267
rect 904 255 944 259
rect -344 188 -340 228
rect -336 188 -332 228
rect -292 188 -288 228
rect -284 188 -280 228
rect -240 188 -236 228
rect -232 188 -228 228
rect -188 188 -184 228
rect -180 188 -176 228
rect -143 196 -139 236
rect -135 196 -131 236
rect -111 196 -107 236
rect -103 196 -99 236
rect 1041 233 1045 273
rect 1049 233 1053 273
rect 1142 234 1146 274
rect 1150 234 1154 274
rect 1194 234 1198 274
rect 1202 234 1206 274
rect 904 212 944 216
rect 904 204 944 208
rect -344 126 -340 166
rect -336 126 -332 166
rect -292 126 -288 166
rect -284 126 -280 166
rect 143 108 147 148
rect 151 108 155 148
rect 181 108 185 148
rect 189 108 193 148
rect 414 116 418 156
rect 422 116 426 156
rect 452 116 456 156
rect 460 116 464 156
rect 378 71 382 91
rect 386 71 390 91
rect 1141 96 1145 136
rect 1149 96 1153 136
rect 1193 96 1197 136
rect 1201 96 1205 136
rect 1245 96 1249 136
rect 1253 96 1257 136
rect 1297 96 1301 136
rect 1305 96 1309 136
rect 1342 104 1346 144
rect 1350 104 1354 144
rect 1374 104 1378 144
rect 1382 104 1386 144
rect 1412 104 1416 124
rect 1420 104 1424 124
rect 904 82 944 86
rect 904 74 944 78
rect 1041 52 1045 92
rect 1049 52 1053 92
rect 904 31 944 35
rect 1141 34 1145 74
rect 1149 34 1153 74
rect 1193 34 1197 74
rect 1201 34 1205 74
rect -345 -23 -341 17
rect -337 -23 -333 17
rect -293 -23 -289 17
rect -285 -23 -281 17
rect -241 -23 -237 17
rect -233 -23 -229 17
rect -189 -23 -185 17
rect -181 -23 -177 17
rect -144 -15 -140 25
rect -136 -15 -132 25
rect -112 -15 -108 25
rect -104 -15 -100 25
rect 6 18 46 22
rect 6 10 46 14
rect 143 -12 147 28
rect 151 -12 155 28
rect 6 -33 46 -29
rect 308 -12 312 28
rect 316 -12 320 28
rect 346 -12 350 28
rect 354 -12 358 28
rect 904 23 944 27
rect -345 -85 -341 -45
rect -337 -85 -333 -45
rect -293 -85 -289 -45
rect -285 -85 -281 -45
rect 6 -41 46 -37
rect 272 -57 276 -37
rect 280 -57 284 -37
rect -353 -227 -349 -187
rect -345 -227 -341 -187
rect -301 -227 -297 -187
rect -293 -227 -289 -187
rect -249 -227 -245 -187
rect -241 -227 -237 -187
rect -197 -227 -193 -187
rect -189 -227 -185 -187
rect -152 -219 -148 -179
rect -144 -219 -140 -179
rect -120 -219 -116 -179
rect -112 -219 -108 -179
rect 143 -182 147 -142
rect 151 -182 155 -142
rect 181 -182 185 -142
rect 189 -182 193 -142
rect 491 -174 495 -134
rect 499 -174 503 -134
rect 529 -174 533 -134
rect 537 -174 541 -134
rect 455 -219 459 -199
rect 463 -219 467 -199
rect -353 -289 -349 -249
rect -345 -289 -341 -249
rect -301 -289 -297 -249
rect -293 -289 -289 -249
rect 6 -272 46 -268
rect 6 -280 46 -276
rect 143 -302 147 -262
rect 151 -302 155 -262
rect 6 -323 46 -319
rect 388 -302 392 -262
rect 396 -302 400 -262
rect 426 -302 430 -262
rect 434 -302 438 -262
rect 6 -331 46 -327
rect 611 -296 615 -256
rect 619 -296 623 -256
rect 649 -296 653 -256
rect 657 -296 661 -256
rect 1140 -303 1144 -263
rect 1148 -303 1152 -263
rect 1192 -303 1196 -263
rect 1200 -303 1204 -263
rect 1244 -303 1248 -263
rect 1252 -303 1256 -263
rect 1296 -303 1300 -263
rect 1304 -303 1308 -263
rect 1341 -295 1345 -255
rect 1349 -295 1353 -255
rect 1373 -295 1377 -255
rect 1381 -295 1385 -255
rect 1411 -295 1415 -275
rect 1419 -295 1423 -275
rect 352 -347 356 -327
rect 360 -347 364 -327
rect 575 -341 579 -321
rect 583 -341 587 -321
rect 904 -330 944 -326
rect 904 -338 944 -334
rect 1041 -360 1045 -320
rect 1049 -360 1053 -320
rect 904 -381 944 -377
rect 1140 -365 1144 -325
rect 1148 -365 1152 -325
rect 1192 -365 1196 -325
rect 1200 -365 1204 -325
rect -354 -438 -350 -398
rect -346 -438 -342 -398
rect -302 -438 -298 -398
rect -294 -438 -290 -398
rect -250 -438 -246 -398
rect -242 -438 -238 -398
rect -198 -438 -194 -398
rect -190 -438 -186 -398
rect -153 -430 -149 -390
rect -145 -430 -141 -390
rect -121 -430 -117 -390
rect -113 -430 -109 -390
rect 316 -428 320 -388
rect 324 -428 328 -388
rect 354 -428 358 -388
rect 362 -428 366 -388
rect 904 -389 944 -385
rect -354 -500 -350 -460
rect -346 -500 -342 -460
rect -302 -500 -298 -460
rect -294 -500 -290 -460
rect 280 -473 284 -453
rect 288 -473 292 -453
rect 445 -458 449 -418
rect 453 -458 457 -418
rect 483 -458 487 -418
rect 491 -458 495 -418
rect 409 -503 413 -483
rect 417 -503 421 -483
rect -359 -633 -355 -593
rect -351 -633 -347 -593
rect -307 -633 -303 -593
rect -299 -633 -295 -593
rect -255 -633 -251 -593
rect -247 -633 -243 -593
rect -203 -633 -199 -593
rect -195 -633 -191 -593
rect -158 -625 -154 -585
rect -150 -625 -146 -585
rect -126 -625 -122 -585
rect -118 -625 -114 -585
rect 143 -599 147 -559
rect 151 -599 155 -559
rect 181 -599 185 -559
rect 189 -599 193 -559
rect 648 -591 652 -551
rect 656 -591 660 -551
rect 686 -591 690 -551
rect 694 -591 698 -551
rect -359 -695 -355 -655
rect -351 -695 -347 -655
rect -307 -695 -303 -655
rect -299 -695 -295 -655
rect 612 -636 616 -616
rect 620 -636 624 -616
rect 6 -689 46 -685
rect 6 -697 46 -693
rect 143 -719 147 -679
rect 151 -719 155 -679
rect 6 -740 46 -736
rect 340 -719 344 -679
rect 348 -719 352 -679
rect 378 -719 382 -679
rect 386 -719 390 -679
rect 6 -748 46 -744
rect 815 -728 819 -688
rect 823 -728 827 -688
rect 853 -728 857 -688
rect 861 -728 865 -688
rect 1140 -717 1144 -677
rect 1148 -717 1152 -677
rect 1192 -717 1196 -677
rect 1200 -717 1204 -677
rect 1244 -717 1248 -677
rect 1252 -717 1256 -677
rect 1296 -717 1300 -677
rect 1304 -717 1308 -677
rect 1341 -709 1345 -669
rect 1349 -709 1353 -669
rect 1373 -709 1377 -669
rect 1381 -709 1385 -669
rect 1411 -709 1415 -689
rect 1419 -709 1423 -689
rect 304 -764 308 -744
rect 312 -764 316 -744
rect 779 -773 783 -753
rect 787 -773 791 -753
rect 905 -762 945 -758
rect 905 -770 945 -766
rect -360 -844 -356 -804
rect -352 -844 -348 -804
rect -308 -844 -304 -804
rect -300 -844 -296 -804
rect -256 -844 -252 -804
rect -248 -844 -244 -804
rect -204 -844 -200 -804
rect -196 -844 -192 -804
rect -159 -836 -155 -796
rect -151 -836 -147 -796
rect -127 -836 -123 -796
rect -119 -836 -115 -796
rect 1042 -792 1046 -752
rect 1050 -792 1054 -752
rect 1140 -779 1144 -739
rect 1148 -779 1152 -739
rect 1192 -779 1196 -739
rect 1200 -779 1204 -739
rect 905 -813 945 -809
rect 905 -821 945 -817
rect -360 -906 -356 -866
rect -352 -906 -348 -866
rect -308 -906 -304 -866
rect -300 -906 -296 -866
rect 340 -863 344 -823
rect 348 -863 352 -823
rect 378 -863 382 -823
rect 386 -863 390 -823
rect 304 -908 308 -888
rect 312 -908 316 -888
rect 469 -893 473 -853
rect 477 -893 481 -853
rect 507 -893 511 -853
rect 515 -893 519 -853
rect 433 -938 437 -918
rect 441 -938 445 -918
rect 644 -947 648 -907
rect 652 -947 656 -907
rect 682 -947 686 -907
rect 690 -947 694 -907
rect 608 -992 612 -972
rect 616 -992 620 -972
rect 343 -1033 347 -993
rect 351 -1033 355 -993
rect 381 -1033 385 -993
rect 389 -1033 393 -993
rect 307 -1078 311 -1058
rect 315 -1078 319 -1058
rect 474 -1063 478 -1023
rect 482 -1063 486 -1023
rect 512 -1063 516 -1023
rect 520 -1063 524 -1023
rect 438 -1108 442 -1088
rect 446 -1108 450 -1088
rect 343 -1177 347 -1137
rect 351 -1177 355 -1137
rect 381 -1177 385 -1137
rect 389 -1177 393 -1137
rect 307 -1222 311 -1202
rect 315 -1222 319 -1202
rect -346 -1335 -342 -1295
rect -338 -1335 -334 -1295
rect -294 -1335 -290 -1295
rect -286 -1335 -282 -1295
rect -242 -1335 -238 -1295
rect -234 -1335 -230 -1295
rect -190 -1335 -186 -1295
rect -182 -1335 -178 -1295
rect -145 -1327 -141 -1287
rect -137 -1327 -133 -1287
rect -113 -1327 -109 -1287
rect -105 -1327 -101 -1287
rect 143 -1300 147 -1260
rect 151 -1300 155 -1260
rect 181 -1300 185 -1260
rect 189 -1300 193 -1260
rect -346 -1397 -342 -1357
rect -338 -1397 -334 -1357
rect -294 -1397 -290 -1357
rect -286 -1397 -282 -1357
rect 6 -1390 46 -1386
rect 6 -1398 46 -1394
rect 143 -1420 147 -1380
rect 151 -1420 155 -1380
rect 6 -1441 46 -1437
rect 352 -1420 356 -1380
rect 360 -1420 364 -1380
rect 390 -1420 394 -1380
rect 398 -1420 402 -1380
rect 506 -1380 510 -1340
rect 514 -1380 518 -1340
rect 544 -1380 548 -1340
rect 552 -1380 556 -1340
rect 6 -1449 46 -1445
rect 470 -1425 474 -1405
rect 478 -1425 482 -1405
rect 1141 -1413 1145 -1373
rect 1149 -1413 1153 -1373
rect 1193 -1413 1197 -1373
rect 1201 -1413 1205 -1373
rect 1245 -1413 1249 -1373
rect 1253 -1413 1257 -1373
rect 1297 -1413 1301 -1373
rect 1305 -1413 1309 -1373
rect 1342 -1405 1346 -1365
rect 1350 -1405 1354 -1365
rect 1374 -1405 1378 -1365
rect 1382 -1405 1386 -1365
rect 1412 -1405 1416 -1385
rect 1420 -1405 1424 -1385
rect 316 -1465 320 -1445
rect 324 -1465 328 -1445
rect 855 -1476 859 -1436
rect 863 -1476 867 -1436
rect 893 -1476 897 -1436
rect 901 -1476 905 -1436
rect 1141 -1475 1145 -1435
rect 1149 -1475 1153 -1435
rect 1193 -1475 1197 -1435
rect 1201 -1475 1205 -1435
rect -347 -1546 -343 -1506
rect -339 -1546 -335 -1506
rect -295 -1546 -291 -1506
rect -287 -1546 -283 -1506
rect -243 -1546 -239 -1506
rect -235 -1546 -231 -1506
rect -191 -1546 -187 -1506
rect -183 -1546 -179 -1506
rect -146 -1538 -142 -1498
rect -138 -1538 -134 -1498
rect -114 -1538 -110 -1498
rect -106 -1538 -102 -1498
rect 819 -1521 823 -1501
rect 827 -1521 831 -1501
rect -347 -1608 -343 -1568
rect -339 -1608 -335 -1568
rect -295 -1608 -291 -1568
rect -287 -1608 -283 -1568
rect 352 -1564 356 -1524
rect 360 -1564 364 -1524
rect 390 -1564 394 -1524
rect 398 -1564 402 -1524
rect 316 -1609 320 -1589
rect 324 -1609 328 -1589
rect 481 -1594 485 -1554
rect 489 -1594 493 -1554
rect 519 -1594 523 -1554
rect 527 -1594 531 -1554
rect 445 -1639 449 -1619
rect 453 -1639 457 -1619
rect 615 -1655 619 -1615
rect 623 -1655 627 -1615
rect 653 -1655 657 -1615
rect 661 -1655 665 -1615
rect 355 -1734 359 -1694
rect 363 -1734 367 -1694
rect 393 -1734 397 -1694
rect 401 -1734 405 -1694
rect 579 -1700 583 -1680
rect 587 -1700 591 -1680
rect 319 -1779 323 -1759
rect 327 -1779 331 -1759
rect 486 -1764 490 -1724
rect 494 -1764 498 -1724
rect 524 -1764 528 -1724
rect 532 -1764 536 -1724
rect 450 -1809 454 -1789
rect 458 -1809 462 -1789
rect 355 -1878 359 -1838
rect 363 -1878 367 -1838
rect 393 -1878 397 -1838
rect 401 -1878 405 -1838
rect 744 -1844 748 -1804
rect 752 -1844 756 -1804
rect 782 -1844 786 -1804
rect 790 -1844 794 -1804
rect 708 -1889 712 -1869
rect 716 -1889 720 -1869
rect 319 -1923 323 -1903
rect 327 -1923 331 -1903
rect 355 -2005 359 -1965
rect 363 -2005 367 -1965
rect 393 -2005 397 -1965
rect 401 -2005 405 -1965
rect 319 -2050 323 -2030
rect 327 -2050 331 -2030
rect 486 -2035 490 -1995
rect 494 -2035 498 -1995
rect 524 -2035 528 -1995
rect 532 -2035 536 -1995
rect 450 -2080 454 -2060
rect 458 -2080 462 -2060
rect 621 -2065 625 -2025
rect 629 -2065 633 -2025
rect 659 -2065 663 -2025
rect 667 -2065 671 -2025
rect 355 -2149 359 -2109
rect 363 -2149 367 -2109
rect 393 -2149 397 -2109
rect 401 -2149 405 -2109
rect 585 -2110 589 -2090
rect 593 -2110 597 -2090
rect 319 -2194 323 -2174
rect 327 -2194 331 -2174
<< psubstratepcontact >>
rect 993 271 997 275
rect 993 247 997 251
rect 993 220 997 224
rect 1405 261 1409 265
rect 1429 261 1433 265
rect 1335 251 1339 255
rect 1359 251 1363 255
rect 1367 251 1371 255
rect 1391 251 1395 255
rect 993 196 997 200
rect 1033 180 1037 184
rect 1057 180 1061 184
rect 1159 180 1163 184
rect 1211 180 1215 184
rect 1263 180 1267 184
rect 1315 180 1319 184
rect -151 143 -147 147
rect -127 143 -123 147
rect -119 143 -115 147
rect -95 143 -91 147
rect -327 72 -323 76
rect -275 72 -271 76
rect -223 72 -219 76
rect -171 72 -167 76
rect 103 62 107 66
rect 993 90 997 94
rect 993 66 997 70
rect 135 55 139 59
rect 159 55 163 59
rect 173 55 177 59
rect 197 55 201 59
rect 406 56 410 60
rect 468 56 472 60
rect 95 26 99 30
rect 993 39 997 43
rect 1404 61 1408 65
rect 1428 61 1432 65
rect 1334 51 1338 55
rect 1358 51 1362 55
rect 1366 51 1370 55
rect 1390 51 1394 55
rect 95 2 99 6
rect 95 -25 99 -21
rect 993 15 997 19
rect 1033 -1 1037 3
rect 1057 -1 1061 3
rect 95 -49 99 -45
rect 1158 -20 1162 -16
rect 1210 -20 1214 -16
rect 1262 -20 1266 -16
rect 1314 -20 1318 -16
rect -152 -68 -148 -64
rect -128 -68 -124 -64
rect -120 -68 -116 -64
rect -96 -68 -92 -64
rect 135 -65 139 -61
rect 159 -65 163 -61
rect 264 -72 268 -68
rect 362 -72 366 -68
rect -328 -139 -324 -135
rect -276 -139 -272 -135
rect -224 -139 -220 -135
rect -172 -139 -168 -135
rect 103 -228 107 -224
rect 135 -235 139 -231
rect 159 -235 163 -231
rect 173 -235 177 -231
rect 197 -235 201 -231
rect 483 -234 487 -230
rect 545 -234 549 -230
rect 95 -264 99 -260
rect -160 -272 -156 -268
rect -136 -272 -132 -268
rect -128 -272 -124 -268
rect -104 -272 -100 -268
rect 95 -288 99 -284
rect 95 -315 99 -311
rect 95 -339 99 -335
rect -336 -343 -332 -339
rect -284 -343 -280 -339
rect -232 -343 -228 -339
rect -180 -343 -176 -339
rect 993 -322 997 -318
rect 135 -355 139 -351
rect 159 -355 163 -351
rect 993 -346 997 -342
rect 603 -356 607 -352
rect 665 -356 669 -352
rect 344 -362 348 -358
rect 442 -362 446 -358
rect 993 -373 997 -369
rect 1403 -338 1407 -334
rect 1427 -338 1431 -334
rect 1333 -348 1337 -344
rect 1357 -348 1361 -344
rect 1365 -348 1369 -344
rect 1389 -348 1393 -344
rect 993 -397 997 -393
rect 1033 -413 1037 -409
rect 1057 -413 1061 -409
rect 1157 -419 1161 -415
rect 1209 -419 1213 -415
rect 1261 -419 1265 -415
rect 1313 -419 1317 -415
rect -161 -483 -157 -479
rect -137 -483 -133 -479
rect -129 -483 -125 -479
rect -105 -483 -101 -479
rect 272 -488 276 -484
rect 370 -488 374 -484
rect 401 -518 405 -514
rect 499 -518 503 -514
rect -337 -554 -333 -550
rect -285 -554 -281 -550
rect -233 -554 -229 -550
rect -181 -554 -177 -550
rect 103 -645 107 -641
rect 135 -652 139 -648
rect 159 -652 163 -648
rect 173 -652 177 -648
rect 197 -652 201 -648
rect 640 -651 644 -647
rect 702 -651 706 -647
rect -166 -678 -162 -674
rect -142 -678 -138 -674
rect -134 -678 -130 -674
rect -110 -678 -106 -674
rect 95 -681 99 -677
rect 95 -705 99 -701
rect 95 -732 99 -728
rect -342 -749 -338 -745
rect -290 -749 -286 -745
rect -238 -749 -234 -745
rect -186 -749 -182 -745
rect 95 -756 99 -752
rect 135 -772 139 -768
rect 159 -772 163 -768
rect 994 -754 998 -750
rect 296 -779 300 -775
rect 394 -779 398 -775
rect 994 -778 998 -774
rect 807 -788 811 -784
rect 869 -788 873 -784
rect 994 -805 998 -801
rect 1403 -752 1407 -748
rect 1427 -752 1431 -748
rect 1333 -762 1337 -758
rect 1357 -762 1361 -758
rect 1365 -762 1369 -758
rect 1389 -762 1393 -758
rect 994 -829 998 -825
rect 1157 -833 1161 -829
rect 1209 -833 1213 -829
rect 1261 -833 1265 -829
rect 1313 -833 1317 -829
rect 1034 -845 1038 -841
rect 1058 -845 1062 -841
rect -167 -889 -163 -885
rect -143 -889 -139 -885
rect -135 -889 -131 -885
rect -111 -889 -107 -885
rect 296 -923 300 -919
rect 394 -923 398 -919
rect 425 -953 429 -949
rect 523 -953 527 -949
rect -343 -960 -339 -956
rect -291 -960 -287 -956
rect -239 -960 -235 -956
rect -187 -960 -183 -956
rect 636 -1007 640 -1003
rect 698 -1007 702 -1003
rect 299 -1093 303 -1089
rect 397 -1093 401 -1089
rect 430 -1123 434 -1119
rect 528 -1123 532 -1119
rect 299 -1237 303 -1233
rect 397 -1237 401 -1233
rect 103 -1346 107 -1342
rect 135 -1353 139 -1349
rect 159 -1353 163 -1349
rect 173 -1353 177 -1349
rect 197 -1353 201 -1349
rect -153 -1380 -149 -1376
rect -129 -1380 -125 -1376
rect -121 -1380 -117 -1376
rect -97 -1380 -93 -1376
rect 95 -1382 99 -1378
rect 95 -1406 99 -1402
rect 95 -1433 99 -1429
rect -329 -1451 -325 -1447
rect -277 -1451 -273 -1447
rect -225 -1451 -221 -1447
rect -173 -1451 -169 -1447
rect 95 -1457 99 -1453
rect 498 -1440 502 -1436
rect 560 -1440 564 -1436
rect 135 -1473 139 -1469
rect 159 -1473 163 -1469
rect 308 -1480 312 -1476
rect 406 -1480 410 -1476
rect 1404 -1448 1408 -1444
rect 1428 -1448 1432 -1444
rect 1334 -1458 1338 -1454
rect 1358 -1458 1362 -1454
rect 1366 -1458 1370 -1454
rect 1390 -1458 1394 -1454
rect 1158 -1529 1162 -1525
rect 1210 -1529 1214 -1525
rect 1262 -1529 1266 -1525
rect 1314 -1529 1318 -1525
rect 847 -1536 851 -1532
rect 909 -1536 913 -1532
rect -154 -1591 -150 -1587
rect -130 -1591 -126 -1587
rect -122 -1591 -118 -1587
rect -98 -1591 -94 -1587
rect 308 -1624 312 -1620
rect 406 -1624 410 -1620
rect 437 -1654 441 -1650
rect 535 -1654 539 -1650
rect -330 -1662 -326 -1658
rect -278 -1662 -274 -1658
rect -226 -1662 -222 -1658
rect -174 -1662 -170 -1658
rect 607 -1715 611 -1711
rect 669 -1715 673 -1711
rect 311 -1794 315 -1790
rect 409 -1794 413 -1790
rect 442 -1824 446 -1820
rect 540 -1824 544 -1820
rect 736 -1904 740 -1900
rect 798 -1904 802 -1900
rect 311 -1938 315 -1934
rect 409 -1938 413 -1934
rect 311 -2065 315 -2061
rect 409 -2065 413 -2061
rect 442 -2095 446 -2091
rect 540 -2095 544 -2091
rect 577 -2125 581 -2121
rect 675 -2125 679 -2121
rect 311 -2209 315 -2205
rect 409 -2209 413 -2205
<< nsubstratencontact >>
rect 1336 352 1340 356
rect 1358 352 1362 356
rect 1368 352 1372 356
rect 1390 352 1394 356
rect 1135 344 1139 348
rect 1157 344 1161 348
rect 1187 344 1191 348
rect 1209 344 1213 348
rect 1239 344 1243 348
rect 1261 344 1265 348
rect 1291 344 1295 348
rect 1313 344 1317 348
rect 1406 332 1410 336
rect 1428 332 1432 336
rect 892 270 896 274
rect 1034 281 1038 285
rect 1056 281 1060 285
rect 892 248 896 252
rect -150 244 -146 248
rect -128 244 -124 248
rect -118 244 -114 248
rect -96 244 -92 248
rect -351 236 -347 240
rect -329 236 -325 240
rect -299 236 -295 240
rect -277 236 -273 240
rect -247 236 -243 240
rect -225 236 -221 240
rect -195 236 -191 240
rect -173 236 -169 240
rect 892 219 896 223
rect 892 197 896 201
rect 407 164 411 168
rect 467 164 471 168
rect 136 156 140 160
rect 158 156 162 160
rect 174 156 178 160
rect 196 156 200 160
rect 1335 152 1339 156
rect 1357 152 1361 156
rect 1367 152 1371 156
rect 1389 152 1393 156
rect 1134 144 1138 148
rect 1156 144 1160 148
rect 1186 144 1190 148
rect 1208 144 1212 148
rect 1238 144 1242 148
rect 1260 144 1264 148
rect 1290 144 1294 148
rect 1312 144 1316 148
rect 892 89 896 93
rect 1034 100 1038 104
rect 1056 100 1060 104
rect 1405 132 1409 136
rect 1427 132 1431 136
rect 892 67 896 71
rect -151 33 -147 37
rect -129 33 -125 37
rect -119 33 -115 37
rect -97 33 -93 37
rect -352 25 -348 29
rect -330 25 -326 29
rect -300 25 -296 29
rect -278 25 -274 29
rect -248 25 -244 29
rect -226 25 -222 29
rect -196 25 -192 29
rect -174 25 -170 29
rect -6 25 -2 29
rect 136 36 140 40
rect 158 36 162 40
rect 301 36 305 40
rect 361 36 365 40
rect 892 38 896 42
rect -6 3 -2 7
rect -6 -26 -2 -22
rect 892 16 896 20
rect -6 -48 -2 -44
rect 484 -126 488 -122
rect 544 -126 548 -122
rect 136 -134 140 -130
rect 158 -134 162 -130
rect 174 -134 178 -130
rect 196 -134 200 -130
rect -159 -171 -155 -167
rect -137 -171 -133 -167
rect -127 -171 -123 -167
rect -105 -171 -101 -167
rect -360 -179 -356 -175
rect -338 -179 -334 -175
rect -308 -179 -304 -175
rect -286 -179 -282 -175
rect -256 -179 -252 -175
rect -234 -179 -230 -175
rect -204 -179 -200 -175
rect -182 -179 -178 -175
rect 604 -248 608 -244
rect 664 -248 668 -244
rect 1334 -247 1338 -243
rect 1356 -247 1360 -243
rect 1366 -247 1370 -243
rect 1388 -247 1392 -243
rect -6 -265 -2 -261
rect 136 -254 140 -250
rect 158 -254 162 -250
rect 381 -254 385 -250
rect 441 -254 445 -250
rect 1133 -255 1137 -251
rect 1155 -255 1159 -251
rect 1185 -255 1189 -251
rect 1207 -255 1211 -251
rect 1237 -255 1241 -251
rect 1259 -255 1263 -251
rect 1289 -255 1293 -251
rect 1311 -255 1315 -251
rect -6 -287 -2 -283
rect -6 -316 -2 -312
rect -6 -338 -2 -334
rect 1404 -267 1408 -263
rect 1426 -267 1430 -263
rect 892 -323 896 -319
rect 1034 -312 1038 -308
rect 1056 -312 1060 -308
rect 892 -345 896 -341
rect 892 -374 896 -370
rect -160 -382 -156 -378
rect -138 -382 -134 -378
rect -128 -382 -124 -378
rect -106 -382 -102 -378
rect 309 -380 313 -376
rect 369 -380 373 -376
rect -361 -390 -357 -386
rect -339 -390 -335 -386
rect -309 -390 -305 -386
rect -287 -390 -283 -386
rect -257 -390 -253 -386
rect -235 -390 -231 -386
rect -205 -390 -201 -386
rect -183 -390 -179 -386
rect 892 -396 896 -392
rect 438 -410 442 -406
rect 498 -410 502 -406
rect 641 -543 645 -539
rect 701 -543 705 -539
rect 136 -551 140 -547
rect 158 -551 162 -547
rect 174 -551 178 -547
rect 196 -551 200 -547
rect -165 -577 -161 -573
rect -143 -577 -139 -573
rect -133 -577 -129 -573
rect -111 -577 -107 -573
rect -366 -585 -362 -581
rect -344 -585 -340 -581
rect -314 -585 -310 -581
rect -292 -585 -288 -581
rect -262 -585 -258 -581
rect -240 -585 -236 -581
rect -210 -585 -206 -581
rect -188 -585 -184 -581
rect 1334 -661 1338 -657
rect 1356 -661 1360 -657
rect 1366 -661 1370 -657
rect 1388 -661 1392 -657
rect -6 -682 -2 -678
rect 136 -671 140 -667
rect 158 -671 162 -667
rect 333 -671 337 -667
rect 393 -671 397 -667
rect 1133 -669 1137 -665
rect 1155 -669 1159 -665
rect 1185 -669 1189 -665
rect 1207 -669 1211 -665
rect 1237 -669 1241 -665
rect 1259 -669 1263 -665
rect 1289 -669 1293 -665
rect 1311 -669 1315 -665
rect -6 -704 -2 -700
rect -6 -733 -2 -729
rect 808 -680 812 -676
rect 868 -680 872 -676
rect -6 -755 -2 -751
rect 1404 -681 1408 -677
rect 1426 -681 1430 -677
rect 893 -755 897 -751
rect 1035 -744 1039 -740
rect 1057 -744 1061 -740
rect -166 -788 -162 -784
rect -144 -788 -140 -784
rect -134 -788 -130 -784
rect -112 -788 -108 -784
rect 893 -777 897 -773
rect -367 -796 -363 -792
rect -345 -796 -341 -792
rect -315 -796 -311 -792
rect -293 -796 -289 -792
rect -263 -796 -259 -792
rect -241 -796 -237 -792
rect -211 -796 -207 -792
rect -189 -796 -185 -792
rect 893 -806 897 -802
rect 333 -815 337 -811
rect 393 -815 397 -811
rect 893 -828 897 -824
rect 462 -845 466 -841
rect 522 -845 526 -841
rect 637 -899 641 -895
rect 697 -899 701 -895
rect 336 -985 340 -981
rect 396 -985 400 -981
rect 467 -1015 471 -1011
rect 527 -1015 531 -1011
rect 336 -1129 340 -1125
rect 396 -1129 400 -1125
rect 136 -1252 140 -1248
rect 158 -1252 162 -1248
rect 174 -1252 178 -1248
rect 196 -1252 200 -1248
rect -152 -1279 -148 -1275
rect -130 -1279 -126 -1275
rect -120 -1279 -116 -1275
rect -98 -1279 -94 -1275
rect -353 -1287 -349 -1283
rect -331 -1287 -327 -1283
rect -301 -1287 -297 -1283
rect -279 -1287 -275 -1283
rect -249 -1287 -245 -1283
rect -227 -1287 -223 -1283
rect -197 -1287 -193 -1283
rect -175 -1287 -171 -1283
rect 499 -1332 503 -1328
rect 559 -1332 563 -1328
rect -6 -1383 -2 -1379
rect 136 -1372 140 -1368
rect 158 -1372 162 -1368
rect 345 -1372 349 -1368
rect 405 -1372 409 -1368
rect -6 -1405 -2 -1401
rect -6 -1434 -2 -1430
rect 1335 -1357 1339 -1353
rect 1357 -1357 1361 -1353
rect 1367 -1357 1371 -1353
rect 1389 -1357 1393 -1353
rect 1134 -1365 1138 -1361
rect 1156 -1365 1160 -1361
rect 1186 -1365 1190 -1361
rect 1208 -1365 1212 -1361
rect 1238 -1365 1242 -1361
rect 1260 -1365 1264 -1361
rect 1290 -1365 1294 -1361
rect 1312 -1365 1316 -1361
rect -6 -1456 -2 -1452
rect 1405 -1377 1409 -1373
rect 1427 -1377 1431 -1373
rect 848 -1428 852 -1424
rect 908 -1428 912 -1424
rect -153 -1490 -149 -1486
rect -131 -1490 -127 -1486
rect -121 -1490 -117 -1486
rect -99 -1490 -95 -1486
rect -354 -1498 -350 -1494
rect -332 -1498 -328 -1494
rect -302 -1498 -298 -1494
rect -280 -1498 -276 -1494
rect -250 -1498 -246 -1494
rect -228 -1498 -224 -1494
rect -198 -1498 -194 -1494
rect -176 -1498 -172 -1494
rect 345 -1516 349 -1512
rect 405 -1516 409 -1512
rect 474 -1546 478 -1542
rect 534 -1546 538 -1542
rect 608 -1607 612 -1603
rect 668 -1607 672 -1603
rect 348 -1686 352 -1682
rect 408 -1686 412 -1682
rect 479 -1716 483 -1712
rect 539 -1716 543 -1712
rect 737 -1796 741 -1792
rect 797 -1796 801 -1792
rect 348 -1830 352 -1826
rect 408 -1830 412 -1826
rect 348 -1957 352 -1953
rect 408 -1957 412 -1953
rect 479 -1987 483 -1983
rect 539 -1987 543 -1983
rect 614 -2017 618 -2013
rect 674 -2017 678 -2013
rect 348 -2101 352 -2097
rect 408 -2101 412 -2097
<< polysilicon >>
rect 1348 344 1350 348
rect 1380 344 1382 348
rect 1147 336 1149 340
rect 1199 336 1201 340
rect 1251 336 1253 340
rect 1303 336 1305 340
rect 1418 324 1420 328
rect 1147 287 1149 296
rect 1199 287 1201 296
rect 1251 287 1253 296
rect 1303 287 1305 296
rect 1014 272 1016 285
rect 1348 284 1350 304
rect 1380 284 1382 304
rect 1418 284 1420 304
rect 1046 273 1048 277
rect 1147 274 1149 278
rect 1199 274 1201 278
rect 900 260 904 262
rect 944 260 964 262
rect 984 260 988 262
rect 1014 248 1016 252
rect -138 236 -136 240
rect -106 236 -104 240
rect 986 242 1016 244
rect 986 239 988 242
rect 1014 240 1016 242
rect -339 228 -337 232
rect -287 228 -285 232
rect -235 228 -233 232
rect -183 228 -181 232
rect 1251 260 1253 269
rect 1303 260 1305 269
rect 1418 270 1420 274
rect 1348 260 1350 264
rect 1380 260 1382 264
rect 1251 237 1253 240
rect 1303 237 1305 240
rect 1014 216 1016 220
rect 1046 213 1048 233
rect 1147 225 1149 234
rect 1199 225 1201 234
rect 1147 213 1149 221
rect 1199 213 1201 221
rect 1251 213 1253 221
rect 1303 213 1305 221
rect 900 209 904 211
rect 944 209 964 211
rect 984 209 988 211
rect -339 179 -337 188
rect -287 179 -285 188
rect -235 179 -233 188
rect -183 179 -181 188
rect -138 176 -136 196
rect -106 176 -104 196
rect 1046 189 1048 193
rect 1147 189 1149 193
rect 1199 189 1201 193
rect 1251 189 1253 193
rect 1303 189 1305 193
rect -339 166 -337 170
rect -287 166 -285 170
rect -235 152 -233 161
rect -183 152 -181 161
rect 419 156 421 160
rect 457 156 459 160
rect -138 152 -136 156
rect -106 152 -104 156
rect 148 148 150 152
rect 186 148 188 152
rect -235 129 -233 132
rect -183 129 -181 132
rect -339 117 -337 126
rect -287 117 -285 126
rect 74 123 118 125
rect 116 121 118 123
rect -339 105 -337 113
rect -287 105 -285 113
rect -235 105 -233 113
rect -183 105 -181 113
rect 383 126 385 130
rect 116 97 118 101
rect 116 89 118 93
rect -339 81 -337 85
rect -287 81 -285 85
rect -235 81 -233 85
rect -183 81 -181 85
rect 148 88 150 108
rect 186 88 188 108
rect 1347 144 1349 148
rect 1379 144 1381 148
rect 1146 136 1148 140
rect 1198 136 1200 140
rect 1250 136 1252 140
rect 1302 136 1304 140
rect 383 91 385 106
rect 419 96 421 116
rect 457 96 459 116
rect 116 53 118 69
rect 1014 91 1016 104
rect 1417 124 1419 128
rect 1046 92 1048 96
rect 900 79 904 81
rect 944 79 964 81
rect 984 79 988 81
rect 419 72 421 76
rect 457 72 459 76
rect 148 64 150 68
rect 186 64 188 68
rect 383 59 385 71
rect 1014 67 1016 71
rect 986 61 1016 63
rect 986 58 988 61
rect 1014 59 1016 61
rect 49 51 118 53
rect -139 25 -137 29
rect -107 25 -105 29
rect 116 27 118 40
rect 1146 87 1148 96
rect 1198 87 1200 96
rect 1250 87 1252 96
rect 1302 87 1304 96
rect 1347 84 1349 104
rect 1379 84 1381 104
rect 1417 84 1419 104
rect 1146 74 1148 78
rect 1198 74 1200 78
rect 1014 35 1016 39
rect 148 28 150 32
rect 313 28 315 32
rect 351 28 353 32
rect 1046 32 1048 52
rect 1250 60 1252 69
rect 1302 60 1304 69
rect 1417 70 1419 74
rect 1347 60 1349 64
rect 1379 60 1381 64
rect 1250 37 1252 40
rect 1302 37 1304 40
rect 900 28 904 30
rect 944 28 964 30
rect 984 28 988 30
rect -340 17 -338 21
rect -288 17 -286 21
rect -236 17 -234 21
rect -184 17 -182 21
rect 2 15 6 17
rect 46 15 66 17
rect 86 15 90 17
rect 116 3 118 7
rect 88 -3 118 -1
rect 88 -6 90 -3
rect 116 -5 118 -3
rect -340 -32 -338 -23
rect -288 -32 -286 -23
rect -236 -32 -234 -23
rect -184 -32 -182 -23
rect -139 -35 -137 -15
rect -107 -35 -105 -15
rect 277 -2 279 6
rect 116 -29 118 -25
rect 148 -32 150 -12
rect 1146 25 1148 34
rect 1198 25 1200 34
rect 1146 13 1148 21
rect 1198 13 1200 21
rect 1250 13 1252 21
rect 1302 13 1304 21
rect 1046 8 1048 12
rect 1146 -11 1148 -7
rect 1198 -11 1200 -7
rect 1250 -11 1252 -7
rect 1302 -11 1304 -7
rect -340 -45 -338 -41
rect -288 -45 -286 -41
rect -236 -59 -234 -50
rect -184 -59 -182 -50
rect 2 -36 6 -34
rect 46 -36 66 -34
rect 86 -36 90 -34
rect 277 -37 279 -22
rect 313 -32 315 -12
rect 351 -32 353 -12
rect -139 -59 -137 -55
rect -107 -59 -105 -55
rect 148 -56 150 -52
rect 313 -56 315 -52
rect 351 -56 353 -52
rect 277 -61 279 -57
rect -236 -82 -234 -79
rect -184 -82 -182 -79
rect -340 -94 -338 -85
rect -288 -94 -286 -85
rect -340 -106 -338 -98
rect -288 -106 -286 -98
rect -236 -106 -234 -98
rect -184 -106 -182 -98
rect -340 -130 -338 -126
rect -288 -130 -286 -126
rect -236 -130 -234 -126
rect -184 -130 -182 -126
rect 496 -134 498 -130
rect 534 -134 536 -130
rect 148 -142 150 -138
rect 186 -142 188 -138
rect 74 -167 118 -165
rect 116 -169 118 -167
rect -147 -179 -145 -175
rect -115 -179 -113 -175
rect -348 -187 -346 -183
rect -296 -187 -294 -183
rect -244 -187 -242 -183
rect -192 -187 -190 -183
rect 460 -164 462 -160
rect 116 -193 118 -189
rect 116 -201 118 -197
rect -348 -236 -346 -227
rect -296 -236 -294 -227
rect -244 -236 -242 -227
rect -192 -236 -190 -227
rect -147 -239 -145 -219
rect -115 -239 -113 -219
rect 148 -202 150 -182
rect 186 -202 188 -182
rect 460 -199 462 -184
rect 496 -194 498 -174
rect 534 -194 536 -174
rect 116 -237 118 -221
rect 496 -218 498 -214
rect 534 -218 536 -214
rect 148 -226 150 -222
rect 186 -226 188 -222
rect 460 -231 462 -219
rect 49 -239 118 -237
rect -348 -249 -346 -245
rect -296 -249 -294 -245
rect -244 -263 -242 -254
rect -192 -263 -190 -254
rect -147 -263 -145 -259
rect -115 -263 -113 -259
rect 116 -263 118 -250
rect 616 -256 618 -252
rect 654 -256 656 -252
rect 1346 -255 1348 -251
rect 1378 -255 1380 -251
rect 148 -262 150 -258
rect 393 -262 395 -258
rect 431 -262 433 -258
rect 2 -275 6 -273
rect 46 -275 66 -273
rect 86 -275 90 -273
rect -244 -286 -242 -283
rect -192 -286 -190 -283
rect 116 -287 118 -283
rect -348 -298 -346 -289
rect -296 -298 -294 -289
rect 88 -293 118 -291
rect 88 -296 90 -293
rect 116 -295 118 -293
rect -348 -310 -346 -302
rect -296 -310 -294 -302
rect -244 -310 -242 -302
rect -192 -310 -190 -302
rect 357 -292 359 -284
rect 116 -319 118 -315
rect 148 -322 150 -302
rect 580 -286 582 -282
rect 2 -326 6 -324
rect 46 -326 66 -324
rect 86 -326 90 -324
rect -348 -334 -346 -330
rect -296 -334 -294 -330
rect -244 -334 -242 -330
rect -192 -334 -190 -330
rect 357 -327 359 -312
rect 393 -322 395 -302
rect 431 -322 433 -302
rect 1145 -263 1147 -259
rect 1197 -263 1199 -259
rect 1249 -263 1251 -259
rect 1301 -263 1303 -259
rect 580 -321 582 -306
rect 616 -316 618 -296
rect 654 -316 656 -296
rect 1416 -275 1418 -271
rect 148 -346 150 -342
rect 1014 -321 1016 -308
rect 1145 -312 1147 -303
rect 1197 -312 1199 -303
rect 1249 -312 1251 -303
rect 1301 -312 1303 -303
rect 1346 -315 1348 -295
rect 1378 -315 1380 -295
rect 1416 -315 1418 -295
rect 1046 -320 1048 -316
rect 900 -333 904 -331
rect 944 -333 964 -331
rect 984 -333 988 -331
rect 616 -340 618 -336
rect 654 -340 656 -336
rect 393 -346 395 -342
rect 431 -346 433 -342
rect 357 -351 359 -347
rect 580 -353 582 -341
rect 1014 -345 1016 -341
rect 986 -351 1016 -349
rect 986 -354 988 -351
rect 1014 -353 1016 -351
rect 1145 -325 1147 -321
rect 1197 -325 1199 -321
rect 1014 -377 1016 -373
rect 1046 -380 1048 -360
rect 1249 -339 1251 -330
rect 1301 -339 1303 -330
rect 1416 -329 1418 -325
rect 1346 -339 1348 -335
rect 1378 -339 1380 -335
rect 1249 -362 1251 -359
rect 1301 -362 1303 -359
rect 1145 -374 1147 -365
rect 1197 -374 1199 -365
rect 900 -384 904 -382
rect 944 -384 964 -382
rect 984 -384 988 -382
rect -148 -390 -146 -386
rect -116 -390 -114 -386
rect 321 -388 323 -384
rect 359 -388 361 -384
rect -349 -398 -347 -394
rect -297 -398 -295 -394
rect -245 -398 -243 -394
rect -193 -398 -191 -394
rect 285 -418 287 -410
rect -349 -447 -347 -438
rect -297 -447 -295 -438
rect -245 -447 -243 -438
rect -193 -447 -191 -438
rect -148 -450 -146 -430
rect -116 -450 -114 -430
rect 1145 -386 1147 -378
rect 1197 -386 1199 -378
rect 1249 -386 1251 -378
rect 1301 -386 1303 -378
rect 1046 -404 1048 -400
rect 1145 -410 1147 -406
rect 1197 -410 1199 -406
rect 1249 -410 1251 -406
rect 1301 -410 1303 -406
rect 450 -418 452 -414
rect 488 -418 490 -414
rect -349 -460 -347 -456
rect -297 -460 -295 -456
rect -245 -474 -243 -465
rect -193 -474 -191 -465
rect 285 -453 287 -438
rect 321 -448 323 -428
rect 359 -448 361 -428
rect 414 -448 416 -440
rect -148 -474 -146 -470
rect -116 -474 -114 -470
rect 321 -472 323 -468
rect 359 -472 361 -468
rect 285 -477 287 -473
rect 414 -483 416 -468
rect 450 -478 452 -458
rect 488 -478 490 -458
rect -245 -497 -243 -494
rect -193 -497 -191 -494
rect -349 -509 -347 -500
rect -297 -509 -295 -500
rect 450 -502 452 -498
rect 488 -502 490 -498
rect 414 -507 416 -503
rect -349 -521 -347 -513
rect -297 -521 -295 -513
rect -245 -521 -243 -513
rect -193 -521 -191 -513
rect -349 -545 -347 -541
rect -297 -545 -295 -541
rect -245 -545 -243 -541
rect -193 -545 -191 -541
rect 653 -551 655 -547
rect 691 -551 693 -547
rect 148 -559 150 -555
rect 186 -559 188 -555
rect -153 -585 -151 -581
rect -121 -585 -119 -581
rect 74 -584 118 -582
rect -354 -593 -352 -589
rect -302 -593 -300 -589
rect -250 -593 -248 -589
rect -198 -593 -196 -589
rect 116 -586 118 -584
rect 617 -581 619 -577
rect 116 -610 118 -606
rect 116 -618 118 -614
rect -354 -642 -352 -633
rect -302 -642 -300 -633
rect -250 -642 -248 -633
rect -198 -642 -196 -633
rect -153 -645 -151 -625
rect -121 -645 -119 -625
rect 148 -619 150 -599
rect 186 -619 188 -599
rect 617 -616 619 -601
rect 653 -611 655 -591
rect 691 -611 693 -591
rect -354 -655 -352 -651
rect -302 -655 -300 -651
rect -250 -669 -248 -660
rect -198 -669 -196 -660
rect 116 -654 118 -638
rect 653 -635 655 -631
rect 691 -635 693 -631
rect 148 -643 150 -639
rect 186 -643 188 -639
rect 617 -648 619 -636
rect 49 -656 118 -654
rect -153 -669 -151 -665
rect -121 -669 -119 -665
rect 116 -680 118 -667
rect 1346 -669 1348 -665
rect 1378 -669 1380 -665
rect 148 -679 150 -675
rect 345 -679 347 -675
rect 383 -679 385 -675
rect -250 -692 -248 -689
rect -198 -692 -196 -689
rect 2 -692 6 -690
rect 46 -692 66 -690
rect 86 -692 90 -690
rect -354 -704 -352 -695
rect -302 -704 -300 -695
rect 116 -704 118 -700
rect -354 -716 -352 -708
rect -302 -716 -300 -708
rect -250 -716 -248 -708
rect -198 -716 -196 -708
rect 88 -710 118 -708
rect 88 -713 90 -710
rect 116 -712 118 -710
rect 309 -709 311 -701
rect 116 -736 118 -732
rect -354 -740 -352 -736
rect -302 -740 -300 -736
rect -250 -740 -248 -736
rect -198 -740 -196 -736
rect 148 -739 150 -719
rect 1145 -677 1147 -673
rect 1197 -677 1199 -673
rect 1249 -677 1251 -673
rect 1301 -677 1303 -673
rect 820 -688 822 -684
rect 858 -688 860 -684
rect 784 -718 786 -714
rect 2 -743 6 -741
rect 46 -743 66 -741
rect 86 -743 90 -741
rect 309 -744 311 -729
rect 345 -739 347 -719
rect 383 -739 385 -719
rect 1416 -689 1418 -685
rect 1145 -726 1147 -717
rect 1197 -726 1199 -717
rect 1249 -726 1251 -717
rect 1301 -726 1303 -717
rect 148 -763 150 -759
rect 784 -753 786 -738
rect 820 -748 822 -728
rect 858 -748 860 -728
rect 1346 -729 1348 -709
rect 1378 -729 1380 -709
rect 1416 -729 1418 -709
rect 1145 -739 1147 -735
rect 1197 -739 1199 -735
rect 345 -763 347 -759
rect 383 -763 385 -759
rect 309 -768 311 -764
rect 1015 -753 1017 -740
rect 1047 -752 1049 -748
rect 901 -765 905 -763
rect 945 -765 965 -763
rect 985 -765 989 -763
rect 820 -772 822 -768
rect 858 -772 860 -768
rect 784 -785 786 -773
rect 1015 -777 1017 -773
rect 987 -783 1017 -781
rect 987 -786 989 -783
rect 1015 -785 1017 -783
rect -154 -796 -152 -792
rect -122 -796 -120 -792
rect -355 -804 -353 -800
rect -303 -804 -301 -800
rect -251 -804 -249 -800
rect -199 -804 -197 -800
rect 1249 -753 1251 -744
rect 1301 -753 1303 -744
rect 1416 -743 1418 -739
rect 1346 -753 1348 -749
rect 1378 -753 1380 -749
rect 1249 -776 1251 -773
rect 1301 -776 1303 -773
rect 1145 -788 1147 -779
rect 1197 -788 1199 -779
rect 1015 -809 1017 -805
rect 1047 -812 1049 -792
rect 1145 -800 1147 -792
rect 1197 -800 1199 -792
rect 1249 -800 1251 -792
rect 1301 -800 1303 -792
rect 901 -816 905 -814
rect 945 -816 965 -814
rect 985 -816 989 -814
rect 345 -823 347 -819
rect 383 -823 385 -819
rect -355 -853 -353 -844
rect -303 -853 -301 -844
rect -251 -853 -249 -844
rect -199 -853 -197 -844
rect -154 -856 -152 -836
rect -122 -856 -120 -836
rect 309 -853 311 -845
rect -355 -866 -353 -862
rect -303 -866 -301 -862
rect -251 -880 -249 -871
rect -199 -880 -197 -871
rect 1145 -824 1147 -820
rect 1197 -824 1199 -820
rect 1249 -824 1251 -820
rect 1301 -824 1303 -820
rect 1047 -836 1049 -832
rect 474 -853 476 -849
rect 512 -853 514 -849
rect -154 -880 -152 -876
rect -122 -880 -120 -876
rect 309 -888 311 -873
rect 345 -883 347 -863
rect 383 -883 385 -863
rect 438 -883 440 -875
rect -251 -903 -249 -900
rect -199 -903 -197 -900
rect -355 -915 -353 -906
rect -303 -915 -301 -906
rect 345 -907 347 -903
rect 383 -907 385 -903
rect 309 -912 311 -908
rect 438 -918 440 -903
rect 474 -913 476 -893
rect 512 -913 514 -893
rect 649 -907 651 -903
rect 687 -907 689 -903
rect -355 -927 -353 -919
rect -303 -927 -301 -919
rect -251 -927 -249 -919
rect -199 -927 -197 -919
rect 474 -937 476 -933
rect 512 -937 514 -933
rect 613 -937 615 -933
rect 438 -942 440 -938
rect -355 -951 -353 -947
rect -303 -951 -301 -947
rect -251 -951 -249 -947
rect -199 -951 -197 -947
rect 613 -972 615 -957
rect 649 -967 651 -947
rect 687 -967 689 -947
rect 348 -993 350 -989
rect 386 -993 388 -989
rect 649 -991 651 -987
rect 687 -991 689 -987
rect 312 -1023 314 -1015
rect 613 -1004 615 -992
rect 479 -1023 481 -1019
rect 517 -1023 519 -1019
rect 312 -1058 314 -1043
rect 348 -1053 350 -1033
rect 386 -1053 388 -1033
rect 443 -1053 445 -1045
rect 348 -1077 350 -1073
rect 386 -1077 388 -1073
rect 312 -1082 314 -1078
rect 443 -1088 445 -1073
rect 479 -1083 481 -1063
rect 517 -1083 519 -1063
rect 479 -1107 481 -1103
rect 517 -1107 519 -1103
rect 443 -1112 445 -1108
rect 348 -1137 350 -1133
rect 386 -1137 388 -1133
rect 312 -1167 314 -1159
rect 312 -1202 314 -1187
rect 348 -1197 350 -1177
rect 386 -1197 388 -1177
rect 348 -1221 350 -1217
rect 386 -1221 388 -1217
rect 312 -1226 314 -1222
rect 148 -1260 150 -1256
rect 186 -1260 188 -1256
rect -140 -1287 -138 -1283
rect -108 -1287 -106 -1283
rect 74 -1285 118 -1283
rect -341 -1295 -339 -1291
rect -289 -1295 -287 -1291
rect -237 -1295 -235 -1291
rect -185 -1295 -183 -1291
rect 116 -1287 118 -1285
rect 116 -1311 118 -1307
rect 116 -1319 118 -1315
rect -341 -1344 -339 -1335
rect -289 -1344 -287 -1335
rect -237 -1344 -235 -1335
rect -185 -1344 -183 -1335
rect -140 -1347 -138 -1327
rect -108 -1347 -106 -1327
rect 148 -1320 150 -1300
rect 186 -1320 188 -1300
rect -341 -1357 -339 -1353
rect -289 -1357 -287 -1353
rect -237 -1371 -235 -1362
rect -185 -1371 -183 -1362
rect 116 -1355 118 -1339
rect 511 -1340 513 -1336
rect 549 -1340 551 -1336
rect 148 -1344 150 -1340
rect 186 -1344 188 -1340
rect 49 -1357 118 -1355
rect -140 -1371 -138 -1367
rect -108 -1371 -106 -1367
rect 116 -1381 118 -1368
rect 475 -1370 477 -1366
rect 148 -1380 150 -1376
rect 357 -1380 359 -1376
rect 395 -1380 397 -1376
rect -237 -1394 -235 -1391
rect -185 -1394 -183 -1391
rect 2 -1393 6 -1391
rect 46 -1393 66 -1391
rect 86 -1393 90 -1391
rect -341 -1406 -339 -1397
rect -289 -1406 -287 -1397
rect 116 -1405 118 -1401
rect -341 -1418 -339 -1410
rect -289 -1418 -287 -1410
rect -237 -1418 -235 -1410
rect -185 -1418 -183 -1410
rect 88 -1411 118 -1409
rect 88 -1414 90 -1411
rect 116 -1413 118 -1411
rect 321 -1410 323 -1402
rect 116 -1437 118 -1433
rect -341 -1442 -339 -1438
rect -289 -1442 -287 -1438
rect -237 -1442 -235 -1438
rect -185 -1442 -183 -1438
rect 148 -1440 150 -1420
rect 1347 -1365 1349 -1361
rect 1379 -1365 1381 -1361
rect 1146 -1373 1148 -1369
rect 1198 -1373 1200 -1369
rect 1250 -1373 1252 -1369
rect 1302 -1373 1304 -1369
rect 475 -1405 477 -1390
rect 511 -1400 513 -1380
rect 549 -1400 551 -1380
rect 2 -1444 6 -1442
rect 46 -1444 66 -1442
rect 86 -1444 90 -1442
rect 321 -1445 323 -1430
rect 357 -1440 359 -1420
rect 395 -1440 397 -1420
rect 1417 -1385 1419 -1381
rect 511 -1424 513 -1420
rect 549 -1424 551 -1420
rect 1146 -1422 1148 -1413
rect 1198 -1422 1200 -1413
rect 1250 -1422 1252 -1413
rect 1302 -1422 1304 -1413
rect 475 -1437 477 -1425
rect 1347 -1425 1349 -1405
rect 1379 -1425 1381 -1405
rect 1417 -1425 1419 -1405
rect 860 -1436 862 -1432
rect 898 -1436 900 -1432
rect 1146 -1435 1148 -1431
rect 1198 -1435 1200 -1431
rect 148 -1464 150 -1460
rect 357 -1464 359 -1460
rect 395 -1464 397 -1460
rect 321 -1469 323 -1465
rect 824 -1466 826 -1462
rect 1250 -1449 1252 -1440
rect 1302 -1449 1304 -1440
rect 1417 -1439 1419 -1435
rect 1347 -1449 1349 -1445
rect 1379 -1449 1381 -1445
rect 1250 -1472 1252 -1469
rect 1302 -1472 1304 -1469
rect -141 -1498 -139 -1494
rect -109 -1498 -107 -1494
rect -342 -1506 -340 -1502
rect -290 -1506 -288 -1502
rect -238 -1506 -236 -1502
rect -186 -1506 -184 -1502
rect 824 -1501 826 -1486
rect 860 -1496 862 -1476
rect 898 -1496 900 -1476
rect 1146 -1484 1148 -1475
rect 1198 -1484 1200 -1475
rect 1146 -1496 1148 -1488
rect 1198 -1496 1200 -1488
rect 1250 -1496 1252 -1488
rect 1302 -1496 1304 -1488
rect 357 -1524 359 -1520
rect 395 -1524 397 -1520
rect 860 -1520 862 -1516
rect 898 -1520 900 -1516
rect 1146 -1520 1148 -1516
rect 1198 -1520 1200 -1516
rect 1250 -1520 1252 -1516
rect 1302 -1520 1304 -1516
rect -342 -1555 -340 -1546
rect -290 -1555 -288 -1546
rect -238 -1555 -236 -1546
rect -186 -1555 -184 -1546
rect -141 -1558 -139 -1538
rect -109 -1558 -107 -1538
rect 321 -1554 323 -1546
rect -342 -1568 -340 -1564
rect -290 -1568 -288 -1564
rect -238 -1582 -236 -1573
rect -186 -1582 -184 -1573
rect 824 -1533 826 -1521
rect 486 -1554 488 -1550
rect 524 -1554 526 -1550
rect -141 -1582 -139 -1578
rect -109 -1582 -107 -1578
rect 321 -1589 323 -1574
rect 357 -1584 359 -1564
rect 395 -1584 397 -1564
rect 450 -1584 452 -1576
rect -238 -1605 -236 -1602
rect -186 -1605 -184 -1602
rect -342 -1617 -340 -1608
rect -290 -1617 -288 -1608
rect 357 -1608 359 -1604
rect 395 -1608 397 -1604
rect 321 -1613 323 -1609
rect 450 -1619 452 -1604
rect 486 -1614 488 -1594
rect 524 -1614 526 -1594
rect -342 -1629 -340 -1621
rect -290 -1629 -288 -1621
rect -238 -1629 -236 -1621
rect -186 -1629 -184 -1621
rect 620 -1615 622 -1611
rect 658 -1615 660 -1611
rect 486 -1638 488 -1634
rect 524 -1638 526 -1634
rect 450 -1643 452 -1639
rect 584 -1645 586 -1641
rect -342 -1653 -340 -1649
rect -290 -1653 -288 -1649
rect -238 -1653 -236 -1649
rect -186 -1653 -184 -1649
rect 584 -1680 586 -1665
rect 620 -1675 622 -1655
rect 658 -1675 660 -1655
rect 360 -1694 362 -1690
rect 398 -1694 400 -1690
rect 324 -1724 326 -1716
rect 620 -1699 622 -1695
rect 658 -1699 660 -1695
rect 584 -1712 586 -1700
rect 491 -1724 493 -1720
rect 529 -1724 531 -1720
rect 324 -1759 326 -1744
rect 360 -1754 362 -1734
rect 398 -1754 400 -1734
rect 455 -1754 457 -1746
rect 360 -1778 362 -1774
rect 398 -1778 400 -1774
rect 324 -1783 326 -1779
rect 455 -1789 457 -1774
rect 491 -1784 493 -1764
rect 529 -1784 531 -1764
rect 749 -1804 751 -1800
rect 787 -1804 789 -1800
rect 491 -1808 493 -1804
rect 529 -1808 531 -1804
rect 455 -1813 457 -1809
rect 713 -1834 715 -1830
rect 360 -1838 362 -1834
rect 398 -1838 400 -1834
rect 324 -1868 326 -1860
rect 713 -1869 715 -1854
rect 749 -1864 751 -1844
rect 787 -1864 789 -1844
rect 324 -1903 326 -1888
rect 360 -1898 362 -1878
rect 398 -1898 400 -1878
rect 749 -1888 751 -1884
rect 787 -1888 789 -1884
rect 713 -1901 715 -1889
rect 360 -1922 362 -1918
rect 398 -1922 400 -1918
rect 324 -1927 326 -1923
rect 360 -1965 362 -1961
rect 398 -1965 400 -1961
rect 324 -1995 326 -1987
rect 491 -1995 493 -1991
rect 529 -1995 531 -1991
rect 324 -2030 326 -2015
rect 360 -2025 362 -2005
rect 398 -2025 400 -2005
rect 455 -2025 457 -2017
rect 626 -2025 628 -2021
rect 664 -2025 666 -2021
rect 360 -2049 362 -2045
rect 398 -2049 400 -2045
rect 324 -2054 326 -2050
rect 455 -2060 457 -2045
rect 491 -2055 493 -2035
rect 529 -2055 531 -2035
rect 590 -2055 592 -2047
rect 491 -2079 493 -2075
rect 529 -2079 531 -2075
rect 455 -2084 457 -2080
rect 590 -2090 592 -2075
rect 626 -2085 628 -2065
rect 664 -2085 666 -2065
rect 360 -2109 362 -2105
rect 398 -2109 400 -2105
rect 324 -2139 326 -2131
rect 626 -2109 628 -2105
rect 664 -2109 666 -2105
rect 590 -2114 592 -2110
rect 324 -2174 326 -2159
rect 360 -2169 362 -2149
rect 398 -2169 400 -2149
rect 360 -2193 362 -2189
rect 398 -2193 400 -2189
rect 324 -2198 326 -2194
<< polycontact >>
rect 1142 287 1147 292
rect 1194 287 1199 292
rect 1246 287 1251 292
rect 1298 287 1303 292
rect 1343 287 1348 292
rect 1009 280 1014 285
rect 1375 287 1380 292
rect 1413 287 1418 292
rect 956 262 961 267
rect 981 239 986 244
rect 1246 264 1251 269
rect 1298 264 1303 269
rect 1041 216 1046 221
rect 956 211 961 216
rect 1142 225 1147 230
rect 1194 225 1199 230
rect 1142 216 1147 221
rect 1194 216 1199 221
rect 1246 216 1251 221
rect 1298 216 1303 221
rect -344 179 -339 184
rect -292 179 -287 184
rect -240 179 -235 184
rect -188 179 -183 184
rect -143 179 -138 184
rect -111 179 -106 184
rect -240 156 -235 161
rect -188 156 -183 161
rect -344 117 -339 122
rect -292 117 -287 122
rect 74 118 79 123
rect -344 108 -339 113
rect -292 108 -287 113
rect -240 108 -235 113
rect -188 108 -183 113
rect 143 91 148 96
rect 181 91 186 96
rect 414 99 419 104
rect 452 99 457 104
rect 1009 99 1014 104
rect 956 81 961 86
rect 378 59 383 64
rect 981 58 986 63
rect 49 46 54 51
rect 111 35 116 40
rect 1141 87 1146 92
rect 1193 87 1198 92
rect 1245 87 1250 92
rect 1297 87 1302 92
rect 1342 87 1347 92
rect 1374 87 1379 92
rect 1412 87 1417 92
rect 1041 35 1046 40
rect 956 30 961 35
rect 1245 64 1250 69
rect 1297 64 1302 69
rect 58 17 63 22
rect 83 -6 88 -1
rect -345 -32 -340 -27
rect -293 -32 -288 -27
rect -241 -32 -236 -27
rect -189 -32 -184 -27
rect -144 -32 -139 -27
rect -112 -32 -107 -27
rect 272 1 277 6
rect 143 -29 148 -24
rect 58 -34 63 -29
rect 1141 25 1146 30
rect 1193 25 1198 30
rect 1141 16 1146 21
rect 1193 16 1198 21
rect 1245 16 1250 21
rect 1297 16 1302 21
rect -241 -55 -236 -50
rect -189 -55 -184 -50
rect 308 -29 313 -24
rect 346 -29 351 -24
rect -345 -94 -340 -89
rect -293 -94 -288 -89
rect -345 -103 -340 -98
rect -293 -103 -288 -98
rect -241 -103 -236 -98
rect -189 -103 -184 -98
rect 74 -172 79 -167
rect 143 -199 148 -194
rect -353 -236 -348 -231
rect -301 -236 -296 -231
rect -249 -236 -244 -231
rect -197 -236 -192 -231
rect -152 -236 -147 -231
rect -120 -236 -115 -231
rect 181 -199 186 -194
rect 491 -191 496 -186
rect 529 -191 534 -186
rect 455 -231 460 -226
rect -249 -259 -244 -254
rect -197 -259 -192 -254
rect 49 -244 54 -239
rect 111 -255 116 -250
rect 58 -273 63 -268
rect -353 -298 -348 -293
rect -301 -298 -296 -293
rect 83 -296 88 -291
rect -353 -307 -348 -302
rect -301 -307 -296 -302
rect -249 -307 -244 -302
rect -197 -307 -192 -302
rect 352 -289 357 -284
rect 143 -319 148 -314
rect 58 -324 63 -319
rect 388 -319 393 -314
rect 426 -319 431 -314
rect 611 -313 616 -308
rect 649 -313 654 -308
rect 1009 -313 1014 -308
rect 1140 -312 1145 -307
rect 1192 -312 1197 -307
rect 1244 -312 1249 -307
rect 1296 -312 1301 -307
rect 1341 -312 1346 -307
rect 1373 -312 1378 -307
rect 1411 -312 1416 -307
rect 956 -331 961 -326
rect 575 -353 580 -348
rect 981 -354 986 -349
rect 1041 -377 1046 -372
rect 956 -382 961 -377
rect 1244 -335 1249 -330
rect 1296 -335 1301 -330
rect 1140 -374 1145 -369
rect 1192 -374 1197 -369
rect 280 -415 285 -410
rect -354 -447 -349 -442
rect -302 -447 -297 -442
rect -250 -447 -245 -442
rect -198 -447 -193 -442
rect -153 -447 -148 -442
rect -121 -447 -116 -442
rect 1140 -383 1145 -378
rect 1192 -383 1197 -378
rect 1244 -383 1249 -378
rect 1296 -383 1301 -378
rect -250 -470 -245 -465
rect -198 -470 -193 -465
rect 316 -445 321 -440
rect 354 -445 359 -440
rect 409 -445 414 -440
rect 445 -475 450 -470
rect 483 -475 488 -470
rect -354 -509 -349 -504
rect -302 -509 -297 -504
rect -354 -518 -349 -513
rect -302 -518 -297 -513
rect -250 -518 -245 -513
rect -198 -518 -193 -513
rect 74 -589 79 -584
rect 143 -616 148 -611
rect -359 -642 -354 -637
rect -307 -642 -302 -637
rect -255 -642 -250 -637
rect -203 -642 -198 -637
rect -158 -642 -153 -637
rect -126 -642 -121 -637
rect 181 -616 186 -611
rect 648 -608 653 -603
rect 686 -608 691 -603
rect -255 -665 -250 -660
rect -203 -665 -198 -660
rect 612 -648 617 -643
rect 49 -661 54 -656
rect 111 -672 116 -667
rect 58 -690 63 -685
rect -359 -704 -354 -699
rect -307 -704 -302 -699
rect -359 -713 -354 -708
rect -307 -713 -302 -708
rect -255 -713 -250 -708
rect -203 -713 -198 -708
rect 83 -713 88 -708
rect 304 -706 309 -701
rect 143 -736 148 -731
rect 58 -741 63 -736
rect 340 -736 345 -731
rect 378 -736 383 -731
rect 1140 -726 1145 -721
rect 1192 -726 1197 -721
rect 1244 -726 1249 -721
rect 1296 -726 1301 -721
rect 1341 -726 1346 -721
rect 815 -745 820 -740
rect 853 -745 858 -740
rect 1373 -726 1378 -721
rect 1411 -726 1416 -721
rect 1010 -745 1015 -740
rect 957 -763 962 -758
rect 779 -785 784 -780
rect 982 -786 987 -781
rect 1244 -749 1249 -744
rect 1296 -749 1301 -744
rect 1140 -788 1145 -783
rect 1192 -788 1197 -783
rect 1042 -809 1047 -804
rect 957 -814 962 -809
rect 1140 -797 1145 -792
rect 1192 -797 1197 -792
rect 1244 -797 1249 -792
rect 1296 -797 1301 -792
rect -360 -853 -355 -848
rect -308 -853 -303 -848
rect -256 -853 -251 -848
rect -204 -853 -199 -848
rect -159 -853 -154 -848
rect -127 -853 -122 -848
rect 304 -850 309 -845
rect -256 -876 -251 -871
rect -204 -876 -199 -871
rect 340 -880 345 -875
rect 378 -880 383 -875
rect 433 -880 438 -875
rect -360 -915 -355 -910
rect -308 -915 -303 -910
rect 469 -910 474 -905
rect 507 -910 512 -905
rect -360 -924 -355 -919
rect -308 -924 -303 -919
rect -256 -924 -251 -919
rect -204 -924 -199 -919
rect 644 -964 649 -959
rect 682 -964 687 -959
rect 307 -1020 312 -1015
rect 608 -1004 613 -999
rect 343 -1050 348 -1045
rect 381 -1050 386 -1045
rect 438 -1050 443 -1045
rect 474 -1080 479 -1075
rect 512 -1080 517 -1075
rect 307 -1164 312 -1159
rect 343 -1194 348 -1189
rect 381 -1194 386 -1189
rect 74 -1290 79 -1285
rect 143 -1317 148 -1312
rect -346 -1344 -341 -1339
rect -294 -1344 -289 -1339
rect -242 -1344 -237 -1339
rect -190 -1344 -185 -1339
rect -145 -1344 -140 -1339
rect -113 -1344 -108 -1339
rect 181 -1317 186 -1312
rect -242 -1367 -237 -1362
rect -190 -1367 -185 -1362
rect 49 -1362 54 -1357
rect 111 -1373 116 -1368
rect 58 -1391 63 -1386
rect -346 -1406 -341 -1401
rect -294 -1406 -289 -1401
rect -346 -1415 -341 -1410
rect -294 -1415 -289 -1410
rect -242 -1415 -237 -1410
rect -190 -1415 -185 -1410
rect 83 -1414 88 -1409
rect 316 -1407 321 -1402
rect 143 -1437 148 -1432
rect 58 -1442 63 -1437
rect 506 -1397 511 -1392
rect 544 -1397 549 -1392
rect 352 -1437 357 -1432
rect 390 -1437 395 -1432
rect 1141 -1422 1146 -1417
rect 1193 -1422 1198 -1417
rect 1245 -1422 1250 -1417
rect 1297 -1422 1302 -1417
rect 1342 -1422 1347 -1417
rect 470 -1437 475 -1432
rect 1374 -1422 1379 -1417
rect 1412 -1422 1417 -1417
rect 1245 -1445 1250 -1440
rect 1297 -1445 1302 -1440
rect 855 -1493 860 -1488
rect 893 -1493 898 -1488
rect 1141 -1484 1146 -1479
rect 1193 -1484 1198 -1479
rect 1141 -1493 1146 -1488
rect 1193 -1493 1198 -1488
rect 1245 -1493 1250 -1488
rect 1297 -1493 1302 -1488
rect -347 -1555 -342 -1550
rect -295 -1555 -290 -1550
rect -243 -1555 -238 -1550
rect -191 -1555 -186 -1550
rect -146 -1555 -141 -1550
rect -114 -1555 -109 -1550
rect 316 -1551 321 -1546
rect -243 -1578 -238 -1573
rect -191 -1578 -186 -1573
rect 819 -1533 824 -1528
rect 352 -1581 357 -1576
rect 390 -1581 395 -1576
rect 445 -1581 450 -1576
rect -347 -1617 -342 -1612
rect -295 -1617 -290 -1612
rect 481 -1611 486 -1606
rect 519 -1611 524 -1606
rect -347 -1626 -342 -1621
rect -295 -1626 -290 -1621
rect -243 -1626 -238 -1621
rect -191 -1626 -186 -1621
rect 615 -1672 620 -1667
rect 653 -1672 658 -1667
rect 319 -1721 324 -1716
rect 579 -1712 584 -1707
rect 355 -1751 360 -1746
rect 393 -1751 398 -1746
rect 450 -1751 455 -1746
rect 486 -1781 491 -1776
rect 524 -1781 529 -1776
rect 319 -1865 324 -1860
rect 744 -1861 749 -1856
rect 782 -1861 787 -1856
rect 355 -1895 360 -1890
rect 393 -1895 398 -1890
rect 708 -1901 713 -1896
rect 319 -1992 324 -1987
rect 355 -2022 360 -2017
rect 393 -2022 398 -2017
rect 450 -2022 455 -2017
rect 486 -2052 491 -2047
rect 524 -2052 529 -2047
rect 585 -2052 590 -2047
rect 621 -2082 626 -2077
rect 659 -2082 664 -2077
rect 319 -2136 324 -2131
rect 355 -2166 360 -2161
rect 393 -2166 398 -2161
<< metal1 >>
rect -418 363 1100 368
rect 1333 356 1397 359
rect 1333 352 1336 356
rect 1340 352 1358 356
rect 1362 352 1368 356
rect 1372 352 1390 356
rect 1394 352 1397 356
rect 1132 348 1320 351
rect 1333 350 1397 352
rect 1132 344 1135 348
rect 1139 344 1157 348
rect 1161 344 1187 348
rect 1191 344 1209 348
rect 1213 344 1239 348
rect 1243 344 1261 348
rect 1265 344 1291 348
rect 1295 344 1313 348
rect 1317 344 1320 348
rect 1132 342 1320 344
rect 1343 344 1347 350
rect 1375 344 1379 350
rect 1142 336 1146 342
rect 1194 336 1198 342
rect 1246 336 1250 342
rect 1298 336 1302 342
rect 1403 336 1435 339
rect 1403 332 1406 336
rect 1410 332 1428 336
rect 1432 332 1435 336
rect 1403 330 1435 332
rect 1413 324 1417 330
rect 1031 285 1063 288
rect 225 280 1009 285
rect 1031 281 1034 285
rect 1038 281 1056 285
rect 1060 281 1063 285
rect 889 274 898 277
rect 889 270 892 274
rect 896 270 898 274
rect 889 267 898 270
rect 956 267 961 280
rect 1031 279 1063 281
rect 1119 287 1142 292
rect 991 275 999 277
rect 991 271 993 275
rect 997 271 999 275
rect 1041 273 1045 279
rect 991 267 999 271
rect 889 263 904 267
rect 889 252 898 263
rect 984 263 999 267
rect 944 255 964 259
rect -153 248 -89 251
rect -153 244 -150 248
rect -146 244 -128 248
rect -124 244 -118 248
rect -114 244 -96 248
rect -92 244 -89 248
rect 889 248 892 252
rect 896 248 898 252
rect 889 245 898 248
rect -354 240 -166 243
rect -153 242 -89 244
rect 956 244 961 255
rect 991 251 999 263
rect 991 247 993 251
rect 997 247 999 251
rect 1009 250 1013 252
rect 991 245 999 247
rect 1002 246 1013 250
rect 1017 248 1021 252
rect -354 236 -351 240
rect -347 236 -329 240
rect -325 236 -299 240
rect -295 236 -277 240
rect -273 236 -247 240
rect -243 236 -225 240
rect -221 236 -195 240
rect -191 236 -173 240
rect -169 236 -166 240
rect -354 234 -166 236
rect -143 236 -139 242
rect -111 236 -107 242
rect 956 239 981 244
rect -344 228 -340 234
rect -292 228 -288 234
rect -240 228 -236 234
rect -188 228 -184 234
rect 1002 235 1006 246
rect 1017 243 1030 248
rect 1017 240 1021 243
rect 234 230 1006 235
rect -367 179 -344 184
rect -367 113 -362 179
rect -336 175 -332 188
rect -344 171 -332 175
rect -314 179 -292 184
rect -344 166 -340 171
rect -349 117 -344 122
rect -336 113 -332 126
rect -314 113 -309 179
rect -284 175 -280 188
rect -232 184 -228 188
rect -180 184 -176 188
rect -135 184 -131 196
rect -103 184 -99 196
rect 889 223 898 226
rect 889 219 892 223
rect 896 219 898 223
rect 889 216 898 219
rect 956 216 961 230
rect 991 224 999 226
rect 991 220 993 224
rect 997 220 999 224
rect 991 216 999 220
rect 889 212 904 216
rect 889 201 898 212
rect 984 212 999 216
rect 944 204 964 208
rect 889 197 892 201
rect 896 197 898 201
rect 889 194 898 197
rect 956 189 961 204
rect 991 200 999 212
rect 991 196 993 200
rect 997 196 999 200
rect 991 194 999 196
rect 1025 221 1030 243
rect 1049 221 1053 233
rect 1119 221 1124 287
rect 1150 283 1154 296
rect 1142 279 1154 283
rect 1172 287 1194 292
rect 1142 274 1146 279
rect 1137 225 1142 230
rect 1150 221 1154 234
rect 1172 221 1177 287
rect 1202 283 1206 296
rect 1254 292 1258 296
rect 1306 292 1310 296
rect 1351 292 1355 304
rect 1383 292 1387 304
rect 1421 292 1425 304
rect 1194 279 1206 283
rect 1224 287 1246 292
rect 1254 287 1298 292
rect 1306 287 1343 292
rect 1351 287 1375 292
rect 1383 287 1413 292
rect 1421 287 1435 292
rect 1194 274 1198 279
rect 1189 225 1194 230
rect 1202 221 1206 234
rect 1224 221 1229 287
rect 1243 264 1246 269
rect 1254 260 1258 287
rect 1246 229 1250 240
rect 1246 225 1258 229
rect 1009 189 1013 220
rect 1025 216 1041 221
rect 1049 216 1142 221
rect 1150 216 1194 221
rect 1202 216 1246 221
rect 1049 213 1053 216
rect 1150 213 1154 216
rect 1202 213 1206 216
rect 1254 213 1258 225
rect 1276 221 1281 287
rect 1295 264 1298 269
rect 1306 260 1310 287
rect 1351 284 1355 287
rect 1383 284 1387 287
rect 1421 284 1425 287
rect 1413 267 1417 274
rect 1403 265 1435 267
rect 1343 257 1347 264
rect 1375 257 1379 264
rect 1403 261 1405 265
rect 1409 261 1429 265
rect 1433 261 1435 265
rect 1403 259 1435 261
rect 1333 255 1397 257
rect 1333 251 1335 255
rect 1339 251 1359 255
rect 1363 251 1367 255
rect 1371 251 1391 255
rect 1395 251 1397 255
rect 1333 249 1397 251
rect 1298 229 1302 240
rect 1298 225 1310 229
rect 1276 216 1298 221
rect 1306 213 1310 225
rect 956 184 1013 189
rect 1041 186 1045 193
rect 1031 184 1063 186
rect 1142 185 1146 193
rect 1194 185 1198 193
rect 1246 185 1250 193
rect 1298 185 1302 193
rect -292 171 -280 175
rect -262 179 -240 184
rect -232 179 -188 184
rect -180 179 -143 184
rect -135 179 -111 184
rect -103 179 -75 184
rect -292 166 -288 171
rect -297 117 -292 122
rect -284 113 -280 126
rect -262 113 -257 179
rect -243 156 -240 161
rect -232 152 -228 179
rect -240 121 -236 132
rect -240 117 -228 121
rect -367 108 -344 113
rect -336 108 -292 113
rect -284 108 -240 113
rect -336 105 -332 108
rect -284 105 -280 108
rect -232 105 -228 117
rect -210 113 -205 179
rect -191 156 -188 161
rect -180 152 -176 179
rect -135 176 -131 179
rect -103 176 -99 179
rect -143 149 -139 156
rect -111 149 -107 156
rect -153 147 -89 149
rect -153 143 -151 147
rect -147 143 -127 147
rect -123 143 -119 147
rect -115 143 -95 147
rect -91 143 -89 147
rect -153 141 -89 143
rect -188 121 -184 132
rect -188 117 -176 121
rect -210 108 -188 113
rect -180 105 -176 117
rect -344 77 -340 85
rect -292 77 -288 85
rect -240 77 -236 85
rect -188 77 -184 85
rect -354 76 -166 77
rect -354 72 -327 76
rect -323 72 -275 76
rect -271 72 -223 76
rect -219 72 -171 76
rect -167 72 -166 76
rect -354 71 -166 72
rect -80 74 -75 179
rect 1031 180 1033 184
rect 1037 180 1057 184
rect 1061 180 1063 184
rect 1031 178 1063 180
rect 1132 184 1320 185
rect 1132 180 1159 184
rect 1163 180 1211 184
rect 1215 180 1263 184
rect 1267 180 1315 184
rect 1319 180 1320 184
rect 1132 179 1320 180
rect 378 168 474 171
rect 378 164 407 168
rect 411 164 467 168
rect 471 164 474 168
rect 1105 166 1132 171
rect 1137 166 1184 171
rect 1189 166 1238 171
rect 1243 166 1290 171
rect 133 160 165 163
rect 133 156 136 160
rect 140 156 158 160
rect 162 156 165 160
rect 133 154 165 156
rect 171 160 203 163
rect 171 156 174 160
rect 178 156 196 160
rect 200 156 203 160
rect 171 154 203 156
rect 378 162 474 164
rect 143 148 147 154
rect 181 148 185 154
rect -22 95 58 100
rect -418 58 -354 63
rect -349 58 -302 63
rect -297 58 -248 63
rect -243 58 -196 63
rect -154 37 -90 40
rect -154 33 -151 37
rect -147 33 -129 37
rect -125 33 -119 37
rect -115 33 -97 37
rect -93 33 -90 37
rect -355 29 -167 32
rect -154 31 -90 33
rect -355 25 -352 29
rect -348 25 -330 29
rect -326 25 -300 29
rect -296 25 -278 29
rect -274 25 -248 29
rect -244 25 -226 29
rect -222 25 -196 29
rect -192 25 -174 29
rect -170 25 -167 29
rect -355 23 -167 25
rect -144 25 -140 31
rect -112 25 -108 31
rect -345 17 -341 23
rect -293 17 -289 23
rect -241 17 -237 23
rect -189 17 -185 23
rect -22 -10 -17 95
rect 74 74 79 118
rect 111 100 115 101
rect 95 95 115 100
rect 119 96 123 101
rect 151 96 155 108
rect 189 96 193 108
rect 378 126 382 162
rect 414 156 418 162
rect 452 156 456 162
rect 1332 156 1396 159
rect 1332 152 1335 156
rect 1339 152 1357 156
rect 1361 152 1367 156
rect 1371 152 1389 156
rect 1393 152 1396 156
rect 1131 148 1319 151
rect 1332 150 1396 152
rect 1131 144 1134 148
rect 1138 144 1156 148
rect 1160 144 1186 148
rect 1190 144 1208 148
rect 1212 144 1238 148
rect 1242 144 1260 148
rect 1264 144 1290 148
rect 1294 144 1312 148
rect 1316 144 1319 148
rect 1131 142 1319 144
rect 1342 144 1346 150
rect 1374 144 1378 150
rect 386 104 390 106
rect 422 104 426 116
rect 460 104 464 116
rect 1141 136 1145 142
rect 1193 136 1197 142
rect 1245 136 1249 142
rect 1297 136 1301 142
rect 1031 104 1063 107
rect 386 99 414 104
rect 422 99 452 104
rect 460 99 1009 104
rect 1031 100 1034 104
rect 1038 100 1056 104
rect 1060 100 1063 104
rect 119 91 143 96
rect 151 91 181 96
rect 189 91 238 96
rect 243 91 383 96
rect 386 91 390 99
rect 422 96 426 99
rect 460 96 464 99
rect 119 89 123 91
rect -9 29 0 32
rect -9 25 -6 29
rect -2 25 0 29
rect -9 22 0 25
rect -9 18 6 22
rect -9 7 0 18
rect 49 14 54 46
rect 74 40 79 69
rect 151 88 155 91
rect 189 88 193 91
rect 111 67 115 69
rect 102 66 115 67
rect 102 62 103 66
rect 107 62 115 66
rect 102 61 115 62
rect 889 93 898 96
rect 889 89 892 93
rect 896 89 898 93
rect 889 86 898 89
rect 956 86 961 99
rect 1031 98 1063 100
rect 991 94 999 96
rect 991 90 993 94
rect 997 90 999 94
rect 1041 92 1045 98
rect 1402 136 1434 139
rect 1402 132 1405 136
rect 1409 132 1427 136
rect 1431 132 1434 136
rect 1402 130 1434 132
rect 1412 124 1416 130
rect 991 86 999 90
rect 889 82 904 86
rect 143 61 147 68
rect 181 61 185 68
rect 133 59 165 61
rect 133 55 135 59
rect 139 55 159 59
rect 163 55 165 59
rect 133 53 165 55
rect 171 59 203 61
rect 171 55 173 59
rect 177 55 197 59
rect 201 55 203 59
rect 171 53 203 55
rect 414 62 418 76
rect 452 62 456 76
rect 889 71 898 82
rect 984 82 999 86
rect 944 74 964 78
rect 889 67 892 71
rect 896 67 898 71
rect 889 64 898 67
rect 956 63 961 74
rect 991 70 999 82
rect 991 66 993 70
rect 997 66 999 70
rect 1009 69 1013 71
rect 991 64 999 66
rect 1002 65 1013 69
rect 1017 67 1021 71
rect 133 40 165 43
rect 58 35 111 40
rect 133 36 136 40
rect 140 36 158 40
rect 162 36 165 40
rect 58 22 63 35
rect 133 34 165 36
rect 298 40 368 43
rect 298 36 301 40
rect 305 36 361 40
rect 365 36 368 40
rect 298 34 368 36
rect 93 30 101 32
rect 93 26 95 30
rect 99 26 101 30
rect 143 28 147 34
rect 308 28 312 34
rect 346 28 350 34
rect 93 22 101 26
rect 86 18 101 22
rect 46 10 66 14
rect -9 3 -6 7
rect -2 3 0 7
rect -9 0 0 3
rect 58 -1 63 10
rect 93 6 101 18
rect 93 2 95 6
rect 99 2 101 6
rect 111 5 115 7
rect 93 0 101 2
rect 104 1 115 5
rect 119 3 123 7
rect 58 -6 83 -1
rect 104 -10 108 1
rect 119 -2 132 3
rect 119 -5 123 -2
rect -368 -32 -345 -27
rect -368 -98 -363 -32
rect -337 -36 -333 -23
rect -345 -40 -333 -36
rect -315 -32 -293 -27
rect -345 -45 -341 -40
rect -350 -94 -345 -89
rect -337 -98 -333 -85
rect -315 -98 -310 -32
rect -285 -36 -281 -23
rect -233 -27 -229 -23
rect -181 -27 -177 -23
rect -136 -27 -132 -15
rect -104 -27 -100 -15
rect -35 -15 108 -10
rect -35 -27 -30 -15
rect -293 -40 -281 -36
rect -263 -32 -241 -27
rect -233 -32 -189 -27
rect -181 -32 -144 -27
rect -136 -32 -112 -27
rect -104 -32 -30 -27
rect -9 -22 0 -19
rect -9 -26 -6 -22
rect -2 -26 0 -22
rect -9 -29 0 -26
rect 58 -29 63 -15
rect 93 -21 101 -19
rect 93 -25 95 -21
rect 99 -25 101 -21
rect 93 -29 101 -25
rect -293 -45 -289 -40
rect -298 -94 -293 -89
rect -285 -98 -281 -85
rect -263 -98 -258 -32
rect -244 -55 -241 -50
rect -233 -59 -229 -32
rect -241 -90 -237 -79
rect -241 -94 -229 -90
rect -368 -103 -345 -98
rect -337 -103 -293 -98
rect -285 -103 -241 -98
rect -337 -106 -333 -103
rect -285 -106 -281 -103
rect -233 -106 -229 -94
rect -211 -98 -206 -32
rect -192 -55 -189 -50
rect -181 -59 -177 -32
rect -136 -35 -132 -32
rect -104 -35 -100 -32
rect -9 -33 6 -29
rect -9 -44 0 -33
rect 86 -33 101 -29
rect 46 -41 66 -37
rect -9 -48 -6 -44
rect -2 -48 0 -44
rect -9 -51 0 -48
rect -144 -62 -140 -55
rect -112 -62 -108 -55
rect 58 -56 63 -41
rect 93 -45 101 -33
rect 93 -49 95 -45
rect 99 -49 101 -45
rect 93 -51 101 -49
rect 127 -24 132 -2
rect 234 1 272 6
rect 151 -24 155 -12
rect 272 -24 276 -22
rect 111 -56 115 -25
rect 127 -29 143 -24
rect 151 -29 220 -24
rect 225 -29 276 -24
rect 280 -24 284 -22
rect 316 -24 320 -12
rect 354 -24 358 -12
rect 378 -24 383 59
rect 404 60 474 62
rect 404 56 406 60
rect 410 56 468 60
rect 472 56 474 60
rect 956 58 981 63
rect 404 54 474 56
rect 1002 54 1006 65
rect 1017 62 1030 67
rect 1017 59 1021 62
rect 894 49 1006 54
rect 889 42 898 45
rect 889 38 892 42
rect 896 38 898 42
rect 889 35 898 38
rect 956 35 961 49
rect 991 43 999 45
rect 991 39 993 43
rect 997 39 999 43
rect 991 35 999 39
rect 889 31 904 35
rect 889 20 898 31
rect 984 31 999 35
rect 944 23 964 27
rect 889 16 892 20
rect 896 16 898 20
rect 889 13 898 16
rect 956 8 961 23
rect 991 19 999 31
rect 991 15 993 19
rect 997 15 999 19
rect 991 13 999 15
rect 1025 40 1030 62
rect 1049 40 1053 52
rect 1118 87 1141 92
rect 1118 40 1123 87
rect 1149 83 1153 96
rect 1009 8 1013 39
rect 1025 35 1041 40
rect 1049 35 1123 40
rect 1049 32 1053 35
rect 956 3 1013 8
rect 1118 21 1123 35
rect 1141 79 1153 83
rect 1171 87 1193 92
rect 1141 74 1145 79
rect 1136 25 1141 30
rect 1149 21 1153 34
rect 1171 21 1176 87
rect 1201 83 1205 96
rect 1253 92 1257 96
rect 1305 92 1309 96
rect 1350 92 1354 104
rect 1382 92 1386 104
rect 1420 92 1424 104
rect 1193 79 1205 83
rect 1223 87 1245 92
rect 1253 87 1297 92
rect 1305 87 1342 92
rect 1350 87 1374 92
rect 1382 87 1412 92
rect 1420 87 1434 92
rect 1193 74 1197 79
rect 1188 25 1193 30
rect 1201 21 1205 34
rect 1223 21 1228 87
rect 1242 64 1245 69
rect 1253 60 1257 87
rect 1245 29 1249 40
rect 1245 25 1257 29
rect 1118 16 1141 21
rect 1149 16 1193 21
rect 1201 16 1245 21
rect 1149 13 1153 16
rect 1201 13 1205 16
rect 1253 13 1257 25
rect 1275 21 1280 87
rect 1294 64 1297 69
rect 1305 60 1309 87
rect 1350 84 1354 87
rect 1382 84 1386 87
rect 1420 84 1424 87
rect 1412 67 1416 74
rect 1402 65 1434 67
rect 1342 57 1346 64
rect 1374 57 1378 64
rect 1402 61 1404 65
rect 1408 61 1428 65
rect 1432 61 1434 65
rect 1402 59 1434 61
rect 1332 55 1396 57
rect 1332 51 1334 55
rect 1338 51 1358 55
rect 1362 51 1366 55
rect 1370 51 1390 55
rect 1394 51 1396 55
rect 1332 49 1396 51
rect 1297 29 1301 40
rect 1297 25 1309 29
rect 1275 16 1297 21
rect 1305 13 1309 25
rect 1041 5 1045 12
rect 1031 3 1063 5
rect 1031 -1 1033 3
rect 1037 -1 1057 3
rect 1061 -1 1063 3
rect 1031 -3 1063 -1
rect 1141 -15 1145 -7
rect 1193 -15 1197 -7
rect 1245 -15 1249 -7
rect 1297 -15 1301 -7
rect 1131 -16 1319 -15
rect 1131 -20 1158 -16
rect 1162 -20 1210 -16
rect 1214 -20 1262 -16
rect 1266 -20 1314 -16
rect 1318 -20 1319 -16
rect 1131 -21 1319 -20
rect 280 -29 308 -24
rect 316 -29 346 -24
rect 354 -29 383 -24
rect 151 -32 155 -29
rect 58 -61 115 -56
rect 280 -37 284 -29
rect 316 -32 320 -29
rect 354 -32 358 -29
rect 143 -59 147 -52
rect 1105 -34 1131 -29
rect 1136 -34 1183 -29
rect 1188 -34 1237 -29
rect 1242 -34 1289 -29
rect 133 -61 165 -59
rect -154 -64 -90 -62
rect -154 -68 -152 -64
rect -148 -68 -128 -64
rect -124 -68 -120 -64
rect -116 -68 -96 -64
rect -92 -68 -90 -64
rect 133 -65 135 -61
rect 139 -65 159 -61
rect 163 -65 165 -61
rect 133 -67 165 -65
rect 272 -66 276 -57
rect 308 -66 312 -52
rect 346 -66 350 -52
rect -154 -70 -90 -68
rect 262 -68 368 -66
rect 262 -72 264 -68
rect 268 -72 362 -68
rect 366 -72 368 -68
rect 262 -74 368 -72
rect -189 -90 -185 -79
rect 252 -86 464 -81
rect -189 -94 -177 -90
rect -211 -103 -189 -98
rect -181 -106 -177 -94
rect 455 -122 551 -119
rect 455 -126 484 -122
rect 488 -126 544 -122
rect 548 -126 551 -122
rect -345 -134 -341 -126
rect -293 -134 -289 -126
rect -241 -134 -237 -126
rect -189 -134 -185 -126
rect 133 -130 165 -127
rect 133 -134 136 -130
rect 140 -134 158 -130
rect 162 -134 165 -130
rect -355 -135 -167 -134
rect -355 -139 -328 -135
rect -324 -139 -276 -135
rect -272 -139 -224 -135
rect -220 -139 -172 -135
rect -168 -139 -167 -135
rect 133 -136 165 -134
rect 171 -130 203 -127
rect 171 -134 174 -130
rect 178 -134 196 -130
rect 200 -134 203 -130
rect 171 -136 203 -134
rect 455 -128 551 -126
rect -355 -140 -167 -139
rect 143 -142 147 -136
rect 181 -142 185 -136
rect -418 -153 -355 -148
rect -350 -153 -303 -148
rect -298 -153 -249 -148
rect -244 -153 -197 -148
rect -162 -167 -98 -164
rect -162 -171 -159 -167
rect -155 -171 -137 -167
rect -133 -171 -127 -167
rect -123 -171 -105 -167
rect -101 -171 -98 -167
rect -363 -175 -175 -172
rect -162 -173 -98 -171
rect -363 -179 -360 -175
rect -356 -179 -338 -175
rect -334 -179 -308 -175
rect -304 -179 -286 -175
rect -282 -179 -256 -175
rect -252 -179 -234 -175
rect -230 -179 -204 -175
rect -200 -179 -182 -175
rect -178 -179 -175 -175
rect -363 -181 -175 -179
rect -152 -179 -148 -173
rect -120 -179 -116 -173
rect -353 -187 -349 -181
rect -301 -187 -297 -181
rect -249 -187 -245 -181
rect -197 -187 -193 -181
rect -376 -236 -353 -231
rect -376 -302 -371 -236
rect -345 -240 -341 -227
rect -353 -244 -341 -240
rect -323 -236 -301 -231
rect -353 -249 -349 -244
rect -358 -298 -353 -293
rect -345 -302 -341 -289
rect -323 -302 -318 -236
rect -293 -240 -289 -227
rect -241 -231 -237 -227
rect -189 -231 -185 -227
rect -144 -231 -140 -219
rect -112 -231 -108 -219
rect -22 -195 58 -190
rect -301 -244 -289 -240
rect -271 -236 -249 -231
rect -241 -236 -197 -231
rect -189 -236 -152 -231
rect -144 -236 -120 -231
rect -112 -236 -99 -231
rect -301 -249 -297 -244
rect -306 -298 -301 -293
rect -293 -302 -289 -289
rect -271 -302 -266 -236
rect -252 -259 -249 -254
rect -241 -263 -237 -236
rect -249 -294 -245 -283
rect -249 -298 -237 -294
rect -376 -307 -353 -302
rect -345 -307 -301 -302
rect -293 -307 -249 -302
rect -345 -310 -341 -307
rect -293 -310 -289 -307
rect -241 -310 -237 -298
rect -219 -302 -214 -236
rect -200 -259 -197 -254
rect -189 -263 -185 -236
rect -144 -239 -140 -236
rect -112 -239 -108 -236
rect -152 -266 -148 -259
rect -120 -266 -116 -259
rect -162 -268 -98 -266
rect -162 -272 -160 -268
rect -156 -272 -136 -268
rect -132 -272 -128 -268
rect -124 -272 -104 -268
rect -100 -272 -98 -268
rect -162 -274 -98 -272
rect -197 -294 -193 -283
rect -197 -298 -185 -294
rect -219 -307 -197 -302
rect -189 -310 -185 -298
rect -22 -300 -17 -195
rect 74 -231 79 -172
rect 111 -190 115 -189
rect 95 -195 115 -190
rect 119 -194 123 -189
rect 151 -194 155 -182
rect 189 -194 193 -182
rect 455 -164 459 -128
rect 491 -134 495 -128
rect 529 -134 533 -128
rect 463 -186 467 -184
rect 499 -186 503 -174
rect 537 -186 541 -174
rect 463 -191 491 -186
rect 499 -191 529 -186
rect 537 -191 560 -186
rect 119 -199 143 -194
rect 151 -199 181 -194
rect 189 -199 256 -194
rect 261 -199 460 -194
rect 463 -199 467 -191
rect 499 -194 503 -191
rect 537 -194 541 -191
rect 119 -201 123 -199
rect 151 -202 155 -199
rect 189 -202 193 -199
rect 111 -223 115 -221
rect 102 -224 115 -223
rect 102 -228 103 -224
rect 107 -228 115 -224
rect 102 -229 115 -228
rect 143 -229 147 -222
rect 181 -229 185 -222
rect -9 -261 0 -258
rect -9 -265 -6 -261
rect -2 -265 0 -261
rect -9 -268 0 -265
rect -9 -272 6 -268
rect -9 -283 0 -272
rect 49 -276 54 -244
rect 74 -250 79 -236
rect 133 -231 165 -229
rect 133 -235 135 -231
rect 139 -235 159 -231
rect 163 -235 165 -231
rect 133 -237 165 -235
rect 171 -231 203 -229
rect 171 -235 173 -231
rect 177 -235 197 -231
rect 201 -235 203 -231
rect 171 -237 203 -235
rect 491 -228 495 -214
rect 529 -228 533 -214
rect 133 -250 165 -247
rect 58 -255 111 -250
rect 133 -254 136 -250
rect 140 -254 158 -250
rect 162 -254 165 -250
rect 58 -268 63 -255
rect 133 -256 165 -254
rect 378 -250 448 -247
rect 378 -254 381 -250
rect 385 -254 441 -250
rect 445 -254 448 -250
rect 378 -256 448 -254
rect 93 -260 101 -258
rect 93 -264 95 -260
rect 99 -264 101 -260
rect 143 -262 147 -256
rect 388 -262 392 -256
rect 426 -262 430 -256
rect 93 -268 101 -264
rect 86 -272 101 -268
rect 46 -280 66 -276
rect -9 -287 -6 -283
rect -2 -287 0 -283
rect -9 -290 0 -287
rect 58 -291 63 -280
rect 93 -284 101 -272
rect 93 -288 95 -284
rect 99 -288 101 -284
rect 111 -285 115 -283
rect 93 -290 101 -288
rect 104 -289 115 -285
rect 119 -287 123 -283
rect 58 -296 83 -291
rect 104 -300 108 -289
rect 119 -292 132 -287
rect 119 -295 123 -292
rect -92 -305 108 -300
rect -353 -338 -349 -330
rect -301 -338 -297 -330
rect -249 -338 -245 -330
rect -197 -338 -193 -330
rect -363 -339 -175 -338
rect -363 -343 -336 -339
rect -332 -343 -284 -339
rect -280 -343 -232 -339
rect -228 -343 -180 -339
rect -176 -343 -175 -339
rect -363 -344 -175 -343
rect -418 -357 -363 -352
rect -358 -357 -311 -352
rect -306 -357 -257 -352
rect -252 -357 -205 -352
rect -163 -378 -99 -375
rect -163 -382 -160 -378
rect -156 -382 -138 -378
rect -134 -382 -128 -378
rect -124 -382 -106 -378
rect -102 -382 -99 -378
rect -364 -386 -176 -383
rect -163 -384 -99 -382
rect -364 -390 -361 -386
rect -357 -390 -339 -386
rect -335 -390 -309 -386
rect -305 -390 -287 -386
rect -283 -390 -257 -386
rect -253 -390 -235 -386
rect -231 -390 -205 -386
rect -201 -390 -183 -386
rect -179 -390 -176 -386
rect -364 -392 -176 -390
rect -153 -390 -149 -384
rect -121 -390 -117 -384
rect -354 -398 -350 -392
rect -302 -398 -298 -392
rect -250 -398 -246 -392
rect -198 -398 -194 -392
rect -377 -447 -354 -442
rect -377 -513 -372 -447
rect -346 -451 -342 -438
rect -354 -455 -342 -451
rect -324 -447 -302 -442
rect -354 -460 -350 -455
rect -359 -509 -354 -504
rect -346 -513 -342 -500
rect -324 -513 -319 -447
rect -294 -451 -290 -438
rect -242 -442 -238 -438
rect -190 -442 -186 -438
rect -145 -442 -141 -430
rect -113 -442 -109 -430
rect -92 -442 -87 -305
rect -9 -312 0 -309
rect -9 -316 -6 -312
rect -2 -316 0 -312
rect -9 -319 0 -316
rect 58 -319 63 -305
rect 93 -311 101 -309
rect 93 -315 95 -311
rect 99 -315 101 -311
rect 93 -319 101 -315
rect -9 -323 6 -319
rect -9 -334 0 -323
rect 86 -323 101 -319
rect 46 -331 66 -327
rect -9 -338 -6 -334
rect -2 -338 0 -334
rect -9 -341 0 -338
rect 58 -346 63 -331
rect 93 -335 101 -323
rect 93 -339 95 -335
rect 99 -339 101 -335
rect 93 -341 101 -339
rect 127 -314 132 -292
rect 243 -289 352 -284
rect 151 -314 155 -302
rect 352 -314 356 -312
rect 111 -346 115 -315
rect 127 -319 143 -314
rect 151 -319 247 -314
rect 252 -319 356 -314
rect 360 -314 364 -312
rect 396 -314 400 -302
rect 434 -314 438 -302
rect 455 -314 460 -231
rect 481 -230 551 -228
rect 481 -234 483 -230
rect 487 -234 545 -230
rect 549 -234 551 -230
rect 481 -236 551 -234
rect 360 -319 388 -314
rect 396 -319 426 -314
rect 434 -319 460 -314
rect 555 -316 560 -191
rect 575 -244 671 -241
rect 575 -248 604 -244
rect 608 -248 664 -244
rect 668 -248 671 -244
rect 1331 -243 1395 -240
rect 1331 -247 1334 -243
rect 1338 -247 1356 -243
rect 1360 -247 1366 -243
rect 1370 -247 1388 -243
rect 1392 -247 1395 -243
rect 575 -250 671 -248
rect 575 -286 579 -250
rect 611 -256 615 -250
rect 649 -256 653 -250
rect 1130 -251 1318 -248
rect 1331 -249 1395 -247
rect 1130 -255 1133 -251
rect 1137 -255 1155 -251
rect 1159 -255 1185 -251
rect 1189 -255 1207 -251
rect 1211 -255 1237 -251
rect 1241 -255 1259 -251
rect 1263 -255 1289 -251
rect 1293 -255 1311 -251
rect 1315 -255 1318 -251
rect 1130 -257 1318 -255
rect 1341 -255 1345 -249
rect 1373 -255 1377 -249
rect 583 -308 587 -306
rect 619 -308 623 -296
rect 657 -308 661 -296
rect 1140 -263 1144 -257
rect 1192 -263 1196 -257
rect 1244 -263 1248 -257
rect 1296 -263 1300 -257
rect 1401 -263 1433 -260
rect 1401 -267 1404 -263
rect 1408 -267 1426 -263
rect 1430 -267 1433 -263
rect 1401 -269 1433 -267
rect 1411 -275 1415 -269
rect 1031 -308 1063 -305
rect 583 -313 611 -308
rect 619 -313 649 -308
rect 657 -313 1009 -308
rect 1031 -312 1034 -308
rect 1038 -312 1056 -308
rect 1060 -312 1063 -308
rect 151 -322 155 -319
rect 58 -351 115 -346
rect 360 -327 364 -319
rect 396 -322 400 -319
rect 434 -322 438 -319
rect 555 -321 580 -316
rect 583 -321 587 -313
rect 619 -316 623 -313
rect 657 -316 661 -313
rect 143 -349 147 -342
rect 889 -319 898 -316
rect 889 -323 892 -319
rect 896 -323 898 -319
rect 889 -326 898 -323
rect 956 -326 961 -313
rect 1031 -314 1063 -312
rect 1117 -312 1140 -307
rect 991 -318 999 -316
rect 991 -322 993 -318
rect 997 -322 999 -318
rect 1041 -320 1045 -314
rect 991 -326 999 -322
rect 889 -330 904 -326
rect 133 -351 165 -349
rect 133 -355 135 -351
rect 139 -355 159 -351
rect 163 -355 165 -351
rect 133 -357 165 -355
rect 352 -356 356 -347
rect 388 -356 392 -342
rect 426 -356 430 -342
rect 565 -353 575 -348
rect 611 -350 615 -336
rect 649 -350 653 -336
rect 889 -341 898 -330
rect 984 -330 999 -326
rect 944 -338 964 -334
rect 889 -345 892 -341
rect 896 -345 898 -341
rect 889 -348 898 -345
rect 956 -349 961 -338
rect 991 -342 999 -330
rect 991 -346 993 -342
rect 997 -346 999 -342
rect 1009 -343 1013 -341
rect 991 -348 999 -346
rect 1002 -347 1013 -343
rect 1017 -345 1021 -341
rect 601 -352 671 -350
rect 342 -358 448 -356
rect 342 -362 344 -358
rect 348 -362 442 -358
rect 446 -362 448 -358
rect 342 -364 448 -362
rect 306 -376 376 -373
rect 306 -380 309 -376
rect 313 -380 369 -376
rect 373 -380 376 -376
rect 306 -382 376 -380
rect 316 -388 320 -382
rect 354 -388 358 -382
rect 225 -415 280 -410
rect 280 -440 284 -438
rect -302 -455 -290 -451
rect -272 -447 -250 -442
rect -242 -447 -198 -442
rect -190 -447 -153 -442
rect -145 -447 -121 -442
rect -113 -447 -87 -442
rect 234 -445 284 -440
rect 435 -406 505 -403
rect 435 -410 438 -406
rect 442 -410 498 -406
rect 502 -410 505 -406
rect 435 -412 505 -410
rect 288 -440 292 -438
rect 324 -440 328 -428
rect 362 -440 366 -428
rect 445 -418 449 -412
rect 483 -418 487 -412
rect 288 -445 316 -440
rect 324 -445 354 -440
rect 362 -445 409 -440
rect -302 -460 -298 -455
rect -307 -509 -302 -504
rect -294 -513 -290 -500
rect -272 -513 -267 -447
rect -253 -470 -250 -465
rect -242 -474 -238 -447
rect -250 -505 -246 -494
rect -250 -509 -238 -505
rect -377 -518 -354 -513
rect -346 -518 -302 -513
rect -294 -518 -250 -513
rect -346 -521 -342 -518
rect -294 -521 -290 -518
rect -242 -521 -238 -509
rect -220 -513 -215 -447
rect -201 -470 -198 -465
rect -190 -474 -186 -447
rect -145 -450 -141 -447
rect -113 -450 -109 -447
rect 288 -453 292 -445
rect 324 -448 328 -445
rect 362 -448 366 -445
rect -153 -477 -149 -470
rect -121 -477 -117 -470
rect -163 -479 -99 -477
rect -163 -483 -161 -479
rect -157 -483 -137 -479
rect -133 -483 -129 -479
rect -125 -483 -105 -479
rect -101 -483 -99 -479
rect 280 -482 284 -473
rect 316 -482 320 -468
rect 354 -482 358 -468
rect 409 -470 413 -468
rect 389 -475 413 -470
rect 417 -470 421 -468
rect 453 -470 457 -458
rect 491 -470 495 -458
rect 565 -470 570 -353
rect 601 -356 603 -352
rect 607 -356 665 -352
rect 669 -356 671 -352
rect 956 -354 981 -349
rect 601 -358 671 -356
rect 1002 -358 1006 -347
rect 1017 -350 1030 -345
rect 1017 -353 1021 -350
rect 894 -363 1006 -358
rect 889 -370 898 -367
rect 889 -374 892 -370
rect 896 -374 898 -370
rect 889 -377 898 -374
rect 956 -377 961 -363
rect 991 -369 999 -367
rect 991 -373 993 -369
rect 997 -373 999 -369
rect 991 -377 999 -373
rect 889 -381 904 -377
rect 889 -392 898 -381
rect 984 -381 999 -377
rect 944 -389 964 -385
rect 889 -396 892 -392
rect 896 -396 898 -392
rect 889 -399 898 -396
rect 956 -404 961 -389
rect 991 -393 999 -381
rect 991 -397 993 -393
rect 997 -397 999 -393
rect 991 -399 999 -397
rect 1025 -372 1030 -350
rect 1049 -372 1053 -360
rect 1117 -372 1122 -312
rect 1148 -316 1152 -303
rect 1140 -320 1152 -316
rect 1170 -312 1192 -307
rect 1140 -325 1144 -320
rect 1009 -404 1013 -373
rect 1025 -377 1041 -372
rect 1049 -377 1122 -372
rect 1135 -374 1140 -369
rect 1049 -380 1053 -377
rect 956 -409 1013 -404
rect 1117 -378 1122 -377
rect 1148 -378 1152 -365
rect 1170 -378 1175 -312
rect 1200 -316 1204 -303
rect 1252 -307 1256 -303
rect 1304 -307 1308 -303
rect 1349 -307 1353 -295
rect 1381 -307 1385 -295
rect 1419 -307 1423 -295
rect 1192 -320 1204 -316
rect 1222 -312 1244 -307
rect 1252 -312 1296 -307
rect 1304 -312 1341 -307
rect 1349 -312 1373 -307
rect 1381 -312 1411 -307
rect 1419 -312 1433 -307
rect 1192 -325 1196 -320
rect 1187 -374 1192 -369
rect 1200 -378 1204 -365
rect 1222 -378 1227 -312
rect 1241 -335 1244 -330
rect 1252 -339 1256 -312
rect 1244 -370 1248 -359
rect 1244 -374 1256 -370
rect 1117 -383 1140 -378
rect 1148 -383 1192 -378
rect 1200 -383 1244 -378
rect 1148 -386 1152 -383
rect 1200 -386 1204 -383
rect 1252 -386 1256 -374
rect 1274 -378 1279 -312
rect 1293 -335 1296 -330
rect 1304 -339 1308 -312
rect 1349 -315 1353 -312
rect 1381 -315 1385 -312
rect 1419 -315 1423 -312
rect 1411 -332 1415 -325
rect 1401 -334 1433 -332
rect 1341 -342 1345 -335
rect 1373 -342 1377 -335
rect 1401 -338 1403 -334
rect 1407 -338 1427 -334
rect 1431 -338 1433 -334
rect 1401 -340 1433 -338
rect 1331 -344 1395 -342
rect 1331 -348 1333 -344
rect 1337 -348 1357 -344
rect 1361 -348 1365 -344
rect 1369 -348 1389 -344
rect 1393 -348 1395 -344
rect 1331 -350 1395 -348
rect 1296 -370 1300 -359
rect 1296 -374 1308 -370
rect 1274 -383 1296 -378
rect 1304 -386 1308 -374
rect 1041 -407 1045 -400
rect 1031 -409 1063 -407
rect 1031 -413 1033 -409
rect 1037 -413 1057 -409
rect 1061 -413 1063 -409
rect 1031 -415 1063 -413
rect 1140 -414 1144 -406
rect 1192 -414 1196 -406
rect 1244 -414 1248 -406
rect 1296 -414 1300 -406
rect 1130 -415 1318 -414
rect 1130 -419 1157 -415
rect 1161 -419 1209 -415
rect 1213 -419 1261 -415
rect 1265 -419 1313 -415
rect 1317 -419 1318 -415
rect 1130 -420 1318 -419
rect 1105 -433 1130 -428
rect 1135 -433 1182 -428
rect 1187 -433 1236 -428
rect 1241 -433 1288 -428
rect 417 -475 445 -470
rect 453 -475 483 -470
rect 491 -475 570 -470
rect -163 -485 -99 -483
rect 270 -484 376 -482
rect 270 -488 272 -484
rect 276 -488 370 -484
rect 374 -488 376 -484
rect 270 -490 376 -488
rect -198 -505 -194 -494
rect 389 -505 395 -475
rect 417 -483 421 -475
rect 453 -478 457 -475
rect 491 -478 495 -475
rect -198 -509 -186 -505
rect -220 -518 -198 -513
rect -190 -521 -186 -509
rect 252 -511 395 -505
rect 409 -512 413 -503
rect 445 -512 449 -498
rect 483 -512 487 -498
rect 399 -514 505 -512
rect 399 -518 401 -514
rect 405 -518 499 -514
rect 503 -518 505 -514
rect 399 -520 505 -518
rect 270 -533 645 -528
rect 612 -539 708 -536
rect -354 -549 -350 -541
rect -302 -549 -298 -541
rect -250 -549 -246 -541
rect -198 -549 -194 -541
rect 612 -543 641 -539
rect 645 -543 701 -539
rect 705 -543 708 -539
rect 133 -547 165 -544
rect -364 -550 -176 -549
rect -364 -554 -337 -550
rect -333 -554 -285 -550
rect -281 -554 -233 -550
rect -229 -554 -181 -550
rect -177 -554 -176 -550
rect 133 -551 136 -547
rect 140 -551 158 -547
rect 162 -551 165 -547
rect 133 -553 165 -551
rect 171 -547 203 -544
rect 171 -551 174 -547
rect 178 -551 196 -547
rect 200 -551 203 -547
rect 171 -553 203 -551
rect 612 -545 708 -543
rect -364 -555 -176 -554
rect 143 -559 147 -553
rect 181 -559 185 -553
rect -418 -568 -364 -563
rect -359 -568 -312 -563
rect -307 -568 -258 -563
rect -253 -568 -206 -563
rect -168 -573 -104 -570
rect -168 -577 -165 -573
rect -161 -577 -143 -573
rect -139 -577 -133 -573
rect -129 -577 -111 -573
rect -107 -577 -104 -573
rect -369 -581 -181 -578
rect -168 -579 -104 -577
rect -369 -585 -366 -581
rect -362 -585 -344 -581
rect -340 -585 -314 -581
rect -310 -585 -292 -581
rect -288 -585 -262 -581
rect -258 -585 -240 -581
rect -236 -585 -210 -581
rect -206 -585 -188 -581
rect -184 -585 -181 -581
rect -369 -587 -181 -585
rect -158 -585 -154 -579
rect -126 -585 -122 -579
rect -359 -593 -355 -587
rect -307 -593 -303 -587
rect -255 -593 -251 -587
rect -203 -593 -199 -587
rect -382 -642 -359 -637
rect -382 -708 -377 -642
rect -351 -646 -347 -633
rect -359 -650 -347 -646
rect -329 -642 -307 -637
rect -359 -655 -355 -650
rect -364 -704 -359 -699
rect -351 -708 -347 -695
rect -329 -708 -324 -642
rect -299 -646 -295 -633
rect -247 -637 -243 -633
rect -195 -637 -191 -633
rect -150 -637 -146 -625
rect -118 -637 -114 -625
rect -22 -612 58 -607
rect -307 -650 -295 -646
rect -277 -642 -255 -637
rect -247 -642 -203 -637
rect -195 -642 -158 -637
rect -150 -642 -126 -637
rect -118 -642 -103 -637
rect -307 -655 -303 -650
rect -312 -704 -307 -699
rect -299 -708 -295 -695
rect -277 -708 -272 -642
rect -258 -665 -255 -660
rect -247 -669 -243 -642
rect -255 -700 -251 -689
rect -255 -704 -243 -700
rect -382 -713 -359 -708
rect -351 -713 -307 -708
rect -299 -713 -255 -708
rect -351 -716 -347 -713
rect -299 -716 -295 -713
rect -247 -716 -243 -704
rect -225 -708 -220 -642
rect -206 -665 -203 -660
rect -195 -669 -191 -642
rect -150 -645 -146 -642
rect -118 -645 -114 -642
rect -158 -672 -154 -665
rect -126 -672 -122 -665
rect -168 -674 -104 -672
rect -168 -678 -166 -674
rect -162 -678 -142 -674
rect -138 -678 -134 -674
rect -130 -678 -110 -674
rect -106 -678 -104 -674
rect -168 -680 -104 -678
rect -203 -700 -199 -689
rect -203 -704 -191 -700
rect -225 -713 -203 -708
rect -195 -716 -191 -704
rect -22 -717 -17 -612
rect 74 -637 79 -589
rect 111 -607 115 -606
rect 95 -612 115 -607
rect 119 -611 123 -606
rect 151 -611 155 -599
rect 189 -611 193 -599
rect 612 -581 616 -545
rect 648 -551 652 -545
rect 686 -551 690 -545
rect 620 -603 624 -601
rect 656 -603 660 -591
rect 694 -603 698 -591
rect 620 -608 648 -603
rect 656 -608 686 -603
rect 694 -608 766 -603
rect 119 -616 143 -611
rect 151 -616 181 -611
rect 189 -616 274 -611
rect 279 -616 617 -611
rect 620 -616 624 -608
rect 656 -611 660 -608
rect 694 -611 698 -608
rect 119 -618 123 -616
rect 151 -619 155 -616
rect 189 -619 193 -616
rect 111 -640 115 -638
rect -9 -678 0 -675
rect -9 -682 -6 -678
rect -2 -682 0 -678
rect -9 -685 0 -682
rect -9 -689 6 -685
rect -9 -700 0 -689
rect 49 -693 54 -661
rect 74 -667 79 -642
rect 102 -641 115 -640
rect 102 -645 103 -641
rect 107 -645 115 -641
rect 102 -646 115 -645
rect 143 -646 147 -639
rect 181 -646 185 -639
rect 133 -648 165 -646
rect 133 -652 135 -648
rect 139 -652 159 -648
rect 163 -652 165 -648
rect 133 -654 165 -652
rect 171 -648 203 -646
rect 171 -652 173 -648
rect 177 -652 197 -648
rect 201 -652 203 -648
rect 171 -654 203 -652
rect 602 -648 612 -643
rect 648 -645 652 -631
rect 686 -645 690 -631
rect 638 -647 708 -645
rect 133 -667 165 -664
rect 58 -672 111 -667
rect 133 -671 136 -667
rect 140 -671 158 -667
rect 162 -671 165 -667
rect 58 -685 63 -672
rect 133 -673 165 -671
rect 330 -667 400 -664
rect 330 -671 333 -667
rect 337 -671 393 -667
rect 397 -671 400 -667
rect 330 -673 400 -671
rect 93 -677 101 -675
rect 93 -681 95 -677
rect 99 -681 101 -677
rect 143 -679 147 -673
rect 340 -679 344 -673
rect 378 -679 382 -673
rect 93 -685 101 -681
rect 86 -689 101 -685
rect 46 -697 66 -693
rect -9 -704 -6 -700
rect -2 -704 0 -700
rect -9 -707 0 -704
rect 58 -708 63 -697
rect 93 -701 101 -689
rect 93 -705 95 -701
rect 99 -705 101 -701
rect 111 -702 115 -700
rect 93 -707 101 -705
rect 104 -706 115 -702
rect 119 -704 123 -700
rect 58 -713 83 -708
rect 104 -717 108 -706
rect 119 -709 132 -704
rect 119 -712 123 -709
rect -96 -722 108 -717
rect -359 -744 -355 -736
rect -307 -744 -303 -736
rect -255 -744 -251 -736
rect -203 -744 -199 -736
rect -369 -745 -181 -744
rect -369 -749 -342 -745
rect -338 -749 -290 -745
rect -286 -749 -238 -745
rect -234 -749 -186 -745
rect -182 -749 -181 -745
rect -369 -750 -181 -749
rect -418 -763 -369 -758
rect -364 -763 -317 -758
rect -312 -763 -263 -758
rect -258 -763 -211 -758
rect -169 -784 -105 -781
rect -169 -788 -166 -784
rect -162 -788 -144 -784
rect -140 -788 -134 -784
rect -130 -788 -112 -784
rect -108 -788 -105 -784
rect -370 -792 -182 -789
rect -169 -790 -105 -788
rect -370 -796 -367 -792
rect -363 -796 -345 -792
rect -341 -796 -315 -792
rect -311 -796 -293 -792
rect -289 -796 -263 -792
rect -259 -796 -241 -792
rect -237 -796 -211 -792
rect -207 -796 -189 -792
rect -185 -796 -182 -792
rect -370 -798 -182 -796
rect -159 -796 -155 -790
rect -127 -796 -123 -790
rect -360 -804 -356 -798
rect -308 -804 -304 -798
rect -256 -804 -252 -798
rect -204 -804 -200 -798
rect -383 -853 -360 -848
rect -383 -919 -378 -853
rect -352 -857 -348 -844
rect -360 -861 -348 -857
rect -330 -853 -308 -848
rect -360 -866 -356 -861
rect -365 -915 -360 -910
rect -352 -919 -348 -906
rect -330 -919 -325 -853
rect -300 -857 -296 -844
rect -248 -848 -244 -844
rect -196 -848 -192 -844
rect -151 -848 -147 -836
rect -119 -848 -115 -836
rect -96 -848 -91 -722
rect -9 -729 0 -726
rect -9 -733 -6 -729
rect -2 -733 0 -729
rect -9 -736 0 -733
rect 58 -736 63 -722
rect 93 -728 101 -726
rect 93 -732 95 -728
rect 99 -732 101 -728
rect 93 -736 101 -732
rect -9 -740 6 -736
rect -9 -751 0 -740
rect 86 -740 101 -736
rect 46 -748 66 -744
rect -9 -755 -6 -751
rect -2 -755 0 -751
rect -9 -758 0 -755
rect 58 -763 63 -748
rect 93 -752 101 -740
rect 93 -756 95 -752
rect 99 -756 101 -752
rect 93 -758 101 -756
rect 127 -731 132 -709
rect 261 -706 304 -701
rect 151 -731 155 -719
rect 304 -731 308 -729
rect 111 -763 115 -732
rect 127 -736 143 -731
rect 151 -736 265 -731
rect 270 -736 308 -731
rect 312 -731 316 -729
rect 348 -731 352 -719
rect 386 -731 390 -719
rect 602 -731 607 -648
rect 638 -651 640 -647
rect 644 -651 702 -647
rect 706 -651 708 -647
rect 638 -653 708 -651
rect 312 -736 340 -731
rect 348 -736 378 -731
rect 386 -736 607 -731
rect 151 -739 155 -736
rect 58 -768 115 -763
rect 312 -744 316 -736
rect 348 -739 352 -736
rect 386 -739 390 -736
rect 143 -766 147 -759
rect 761 -748 766 -608
rect 1331 -657 1395 -654
rect 1331 -661 1334 -657
rect 1338 -661 1356 -657
rect 1360 -661 1366 -657
rect 1370 -661 1388 -657
rect 1392 -661 1395 -657
rect 1130 -665 1318 -662
rect 1331 -663 1395 -661
rect 1130 -669 1133 -665
rect 1137 -669 1155 -665
rect 1159 -669 1185 -665
rect 1189 -669 1207 -665
rect 1211 -669 1237 -665
rect 1241 -669 1259 -665
rect 1263 -669 1289 -665
rect 1293 -669 1311 -665
rect 1315 -669 1318 -665
rect 1130 -671 1318 -669
rect 1341 -669 1345 -663
rect 1373 -669 1377 -663
rect 779 -676 875 -673
rect 779 -680 808 -676
rect 812 -680 868 -676
rect 872 -680 875 -676
rect 779 -682 875 -680
rect 1140 -677 1144 -671
rect 1192 -677 1196 -671
rect 1244 -677 1248 -671
rect 1296 -677 1300 -671
rect 779 -718 783 -682
rect 815 -688 819 -682
rect 853 -688 857 -682
rect 1401 -677 1433 -674
rect 1401 -681 1404 -677
rect 1408 -681 1426 -677
rect 1430 -681 1433 -677
rect 1401 -683 1433 -681
rect 1411 -689 1415 -683
rect 787 -740 791 -738
rect 823 -740 827 -728
rect 861 -740 865 -728
rect 1117 -726 1140 -721
rect 1032 -740 1064 -737
rect 787 -745 815 -740
rect 823 -745 853 -740
rect 861 -745 1010 -740
rect 1032 -744 1035 -740
rect 1039 -744 1057 -740
rect 1061 -744 1064 -740
rect 761 -753 784 -748
rect 787 -753 791 -745
rect 823 -748 827 -745
rect 861 -748 865 -745
rect 133 -768 165 -766
rect 133 -772 135 -768
rect 139 -772 159 -768
rect 163 -772 165 -768
rect 133 -774 165 -772
rect 304 -773 308 -764
rect 340 -773 344 -759
rect 378 -773 382 -759
rect 890 -751 899 -748
rect 890 -755 893 -751
rect 897 -755 899 -751
rect 890 -758 899 -755
rect 957 -758 962 -745
rect 1032 -746 1064 -744
rect 992 -750 1000 -748
rect 992 -754 994 -750
rect 998 -754 1000 -750
rect 1042 -752 1046 -746
rect 992 -758 1000 -754
rect 890 -762 905 -758
rect 294 -775 400 -773
rect 294 -779 296 -775
rect 300 -779 394 -775
rect 398 -779 400 -775
rect 294 -781 400 -779
rect 761 -785 779 -780
rect 815 -782 819 -768
rect 853 -782 857 -768
rect 890 -773 899 -762
rect 985 -762 1000 -758
rect 945 -770 965 -766
rect 890 -777 893 -773
rect 897 -777 899 -773
rect 890 -780 899 -777
rect 957 -781 962 -770
rect 992 -774 1000 -762
rect 992 -778 994 -774
rect 998 -778 1000 -774
rect 1010 -775 1014 -773
rect 992 -780 1000 -778
rect 1003 -779 1014 -775
rect 1018 -777 1022 -773
rect 805 -784 875 -782
rect 330 -811 400 -808
rect 330 -815 333 -811
rect 337 -815 393 -811
rect 397 -815 400 -811
rect 330 -817 400 -815
rect 340 -823 344 -817
rect 378 -823 382 -817
rect -308 -861 -296 -857
rect -278 -853 -256 -848
rect -248 -853 -204 -848
rect -196 -853 -159 -848
rect -151 -853 -127 -848
rect -119 -853 -91 -848
rect 243 -850 304 -845
rect -308 -866 -304 -861
rect -313 -915 -308 -910
rect -300 -919 -296 -906
rect -278 -919 -273 -853
rect -259 -876 -256 -871
rect -248 -880 -244 -853
rect -256 -911 -252 -900
rect -256 -915 -244 -911
rect -383 -924 -360 -919
rect -352 -924 -308 -919
rect -300 -924 -256 -919
rect -352 -927 -348 -924
rect -300 -927 -296 -924
rect -248 -927 -244 -915
rect -226 -919 -221 -853
rect -207 -876 -204 -871
rect -196 -880 -192 -853
rect -151 -856 -147 -853
rect -119 -856 -115 -853
rect 304 -875 308 -873
rect -159 -883 -155 -876
rect -127 -883 -123 -876
rect 252 -880 308 -875
rect 459 -841 529 -838
rect 459 -845 462 -841
rect 466 -845 522 -841
rect 526 -845 529 -841
rect 459 -847 529 -845
rect 312 -875 316 -873
rect 348 -875 352 -863
rect 386 -875 390 -863
rect 469 -853 473 -847
rect 507 -853 511 -847
rect 312 -880 340 -875
rect 348 -880 378 -875
rect 386 -880 433 -875
rect -169 -885 -105 -883
rect -169 -889 -167 -885
rect -163 -889 -143 -885
rect -139 -889 -135 -885
rect -131 -889 -111 -885
rect -107 -889 -105 -885
rect 312 -888 316 -880
rect 348 -883 352 -880
rect 386 -883 390 -880
rect -169 -891 -105 -889
rect -204 -911 -200 -900
rect -204 -915 -192 -911
rect -226 -924 -204 -919
rect -196 -927 -192 -915
rect 304 -917 308 -908
rect 340 -917 344 -903
rect 378 -917 382 -903
rect 433 -905 437 -903
rect 413 -910 437 -905
rect 441 -905 445 -903
rect 477 -905 481 -893
rect 515 -905 519 -893
rect 608 -895 704 -892
rect 608 -899 637 -895
rect 641 -899 697 -895
rect 701 -899 704 -895
rect 608 -901 704 -899
rect 441 -910 469 -905
rect 477 -910 507 -905
rect 515 -910 581 -905
rect 294 -919 400 -917
rect 294 -923 296 -919
rect 300 -923 394 -919
rect 398 -923 400 -919
rect 294 -925 400 -923
rect 413 -940 419 -910
rect 441 -918 445 -910
rect 477 -913 481 -910
rect 515 -913 519 -910
rect 270 -945 419 -940
rect 433 -947 437 -938
rect 469 -947 473 -933
rect 507 -947 511 -933
rect -360 -955 -356 -947
rect -308 -955 -304 -947
rect -256 -955 -252 -947
rect -204 -955 -200 -947
rect 423 -949 529 -947
rect 423 -953 425 -949
rect 429 -953 523 -949
rect 527 -953 529 -949
rect 423 -955 529 -953
rect -370 -956 -182 -955
rect -370 -960 -343 -956
rect -339 -960 -291 -956
rect -287 -960 -239 -956
rect -235 -960 -187 -956
rect -183 -960 -182 -956
rect -370 -961 -182 -960
rect 576 -967 581 -910
rect 608 -937 612 -901
rect 644 -907 648 -901
rect 682 -907 686 -901
rect 616 -959 620 -957
rect 652 -959 656 -947
rect 690 -959 694 -947
rect 761 -959 766 -785
rect 805 -788 807 -784
rect 811 -788 869 -784
rect 873 -788 875 -784
rect 957 -786 982 -781
rect 805 -790 875 -788
rect 1003 -790 1007 -779
rect 1018 -782 1031 -777
rect 1018 -785 1022 -782
rect 895 -795 1007 -790
rect 890 -802 899 -799
rect 890 -806 893 -802
rect 897 -806 899 -802
rect 890 -809 899 -806
rect 957 -809 962 -795
rect 992 -801 1000 -799
rect 992 -805 994 -801
rect 998 -805 1000 -801
rect 992 -809 1000 -805
rect 890 -813 905 -809
rect 890 -824 899 -813
rect 985 -813 1000 -809
rect 945 -821 965 -817
rect 890 -828 893 -824
rect 897 -828 899 -824
rect 890 -831 899 -828
rect 957 -836 962 -821
rect 992 -825 1000 -813
rect 992 -829 994 -825
rect 998 -829 1000 -825
rect 992 -831 1000 -829
rect 1026 -804 1031 -782
rect 1117 -792 1122 -726
rect 1148 -730 1152 -717
rect 1140 -734 1152 -730
rect 1170 -726 1192 -721
rect 1140 -739 1144 -734
rect 1135 -788 1140 -783
rect 1148 -792 1152 -779
rect 1170 -792 1175 -726
rect 1200 -730 1204 -717
rect 1252 -721 1256 -717
rect 1304 -721 1308 -717
rect 1349 -721 1353 -709
rect 1381 -721 1385 -709
rect 1419 -721 1423 -709
rect 1192 -734 1204 -730
rect 1222 -726 1244 -721
rect 1252 -726 1296 -721
rect 1304 -726 1341 -721
rect 1349 -726 1373 -721
rect 1381 -726 1411 -721
rect 1419 -726 1433 -721
rect 1192 -739 1196 -734
rect 1187 -788 1192 -783
rect 1200 -792 1204 -779
rect 1222 -792 1227 -726
rect 1241 -749 1244 -744
rect 1252 -753 1256 -726
rect 1244 -784 1248 -773
rect 1244 -788 1256 -784
rect 1050 -804 1054 -792
rect 1089 -797 1140 -792
rect 1148 -797 1192 -792
rect 1200 -797 1244 -792
rect 1089 -804 1094 -797
rect 1148 -800 1152 -797
rect 1200 -800 1204 -797
rect 1252 -800 1256 -788
rect 1274 -792 1279 -726
rect 1293 -749 1296 -744
rect 1304 -753 1308 -726
rect 1349 -729 1353 -726
rect 1381 -729 1385 -726
rect 1419 -729 1423 -726
rect 1411 -746 1415 -739
rect 1401 -748 1433 -746
rect 1341 -756 1345 -749
rect 1373 -756 1377 -749
rect 1401 -752 1403 -748
rect 1407 -752 1427 -748
rect 1431 -752 1433 -748
rect 1401 -754 1433 -752
rect 1331 -758 1395 -756
rect 1331 -762 1333 -758
rect 1337 -762 1357 -758
rect 1361 -762 1365 -758
rect 1369 -762 1389 -758
rect 1393 -762 1395 -758
rect 1331 -764 1395 -762
rect 1296 -784 1300 -773
rect 1296 -788 1308 -784
rect 1274 -797 1296 -792
rect 1304 -800 1308 -788
rect 1010 -836 1014 -805
rect 1026 -809 1042 -804
rect 1050 -809 1094 -804
rect 1050 -812 1054 -809
rect 957 -841 1014 -836
rect 1140 -828 1144 -820
rect 1192 -828 1196 -820
rect 1244 -828 1248 -820
rect 1296 -828 1300 -820
rect 1130 -829 1318 -828
rect 1042 -839 1046 -832
rect 1130 -833 1157 -829
rect 1161 -833 1209 -829
rect 1213 -833 1261 -829
rect 1265 -833 1313 -829
rect 1317 -833 1318 -829
rect 1130 -834 1318 -833
rect 1032 -841 1064 -839
rect 1032 -845 1034 -841
rect 1038 -845 1058 -841
rect 1062 -845 1064 -841
rect 1032 -847 1064 -845
rect 1105 -847 1130 -842
rect 1135 -847 1182 -842
rect 1187 -847 1236 -842
rect 1241 -847 1288 -842
rect 616 -964 644 -959
rect 652 -964 682 -959
rect 690 -964 766 -959
rect -418 -974 -370 -969
rect -365 -974 -318 -969
rect -313 -974 -264 -969
rect -259 -974 -212 -969
rect 576 -972 613 -967
rect 616 -972 620 -964
rect 652 -967 656 -964
rect 690 -967 694 -964
rect 333 -981 403 -978
rect 333 -985 336 -981
rect 340 -985 396 -981
rect 400 -985 403 -981
rect 333 -987 403 -985
rect 343 -993 347 -987
rect 381 -993 385 -987
rect 225 -1020 307 -1015
rect 307 -1045 311 -1043
rect 234 -1050 311 -1045
rect 598 -1004 608 -999
rect 644 -1001 648 -987
rect 682 -1001 686 -987
rect 634 -1003 704 -1001
rect 464 -1011 534 -1008
rect 464 -1015 467 -1011
rect 471 -1015 527 -1011
rect 531 -1015 534 -1011
rect 464 -1017 534 -1015
rect 315 -1045 319 -1043
rect 351 -1045 355 -1033
rect 389 -1045 393 -1033
rect 474 -1023 478 -1017
rect 512 -1023 516 -1017
rect 315 -1050 343 -1045
rect 351 -1050 381 -1045
rect 389 -1050 438 -1045
rect 315 -1058 319 -1050
rect 351 -1053 355 -1050
rect 389 -1053 393 -1050
rect 307 -1087 311 -1078
rect 343 -1087 347 -1073
rect 381 -1087 385 -1073
rect 438 -1075 442 -1073
rect 408 -1080 442 -1075
rect 446 -1075 450 -1073
rect 482 -1075 486 -1063
rect 520 -1075 524 -1063
rect 598 -1075 604 -1004
rect 634 -1007 636 -1003
rect 640 -1007 698 -1003
rect 702 -1007 704 -1003
rect 634 -1009 704 -1007
rect 446 -1080 474 -1075
rect 482 -1080 512 -1075
rect 520 -1080 604 -1075
rect 297 -1089 403 -1087
rect 297 -1093 299 -1089
rect 303 -1093 397 -1089
rect 401 -1093 403 -1089
rect 297 -1095 403 -1093
rect 333 -1125 403 -1122
rect 333 -1129 336 -1125
rect 340 -1129 396 -1125
rect 400 -1129 403 -1125
rect 333 -1131 403 -1129
rect 343 -1137 347 -1131
rect 381 -1137 385 -1131
rect 252 -1164 307 -1159
rect 307 -1189 311 -1187
rect 270 -1194 311 -1189
rect 315 -1189 319 -1187
rect 351 -1189 355 -1177
rect 389 -1189 393 -1177
rect 408 -1189 413 -1080
rect 446 -1088 450 -1080
rect 482 -1083 486 -1080
rect 520 -1083 524 -1080
rect 438 -1117 442 -1108
rect 474 -1117 478 -1103
rect 512 -1117 516 -1103
rect 428 -1119 534 -1117
rect 428 -1123 430 -1119
rect 434 -1123 528 -1119
rect 532 -1123 534 -1119
rect 428 -1125 534 -1123
rect 315 -1194 343 -1189
rect 351 -1194 381 -1189
rect 389 -1194 413 -1189
rect 315 -1202 319 -1194
rect 351 -1197 355 -1194
rect 389 -1197 393 -1194
rect 307 -1231 311 -1222
rect 343 -1231 347 -1217
rect 381 -1231 385 -1217
rect 297 -1233 403 -1231
rect 297 -1237 299 -1233
rect 303 -1237 397 -1233
rect 401 -1237 403 -1233
rect 297 -1239 403 -1237
rect 133 -1248 165 -1245
rect 133 -1252 136 -1248
rect 140 -1252 158 -1248
rect 162 -1252 165 -1248
rect 133 -1254 165 -1252
rect 171 -1248 203 -1245
rect 171 -1252 174 -1248
rect 178 -1252 196 -1248
rect 200 -1252 203 -1248
rect 288 -1249 853 -1244
rect 171 -1254 203 -1252
rect 143 -1260 147 -1254
rect 181 -1260 185 -1254
rect -155 -1275 -91 -1272
rect -155 -1279 -152 -1275
rect -148 -1279 -130 -1275
rect -126 -1279 -120 -1275
rect -116 -1279 -98 -1275
rect -94 -1279 -91 -1275
rect -356 -1283 -168 -1280
rect -155 -1281 -91 -1279
rect -356 -1287 -353 -1283
rect -349 -1287 -331 -1283
rect -327 -1287 -301 -1283
rect -297 -1287 -279 -1283
rect -275 -1287 -249 -1283
rect -245 -1287 -227 -1283
rect -223 -1287 -197 -1283
rect -193 -1287 -175 -1283
rect -171 -1287 -168 -1283
rect -356 -1289 -168 -1287
rect -145 -1287 -141 -1281
rect -113 -1287 -109 -1281
rect -346 -1295 -342 -1289
rect -294 -1295 -290 -1289
rect -242 -1295 -238 -1289
rect -190 -1295 -186 -1289
rect -369 -1344 -346 -1339
rect -369 -1410 -364 -1344
rect -338 -1348 -334 -1335
rect -346 -1352 -334 -1348
rect -316 -1344 -294 -1339
rect -346 -1357 -342 -1352
rect -351 -1406 -346 -1401
rect -338 -1410 -334 -1397
rect -316 -1410 -311 -1344
rect -286 -1348 -282 -1335
rect -234 -1339 -230 -1335
rect -182 -1339 -178 -1335
rect -137 -1339 -133 -1327
rect -105 -1339 -101 -1327
rect -22 -1313 58 -1308
rect -294 -1352 -282 -1348
rect -264 -1344 -242 -1339
rect -234 -1344 -190 -1339
rect -182 -1344 -145 -1339
rect -137 -1344 -113 -1339
rect -105 -1344 -93 -1339
rect -294 -1357 -290 -1352
rect -299 -1406 -294 -1401
rect -286 -1410 -282 -1397
rect -264 -1410 -259 -1344
rect -245 -1367 -242 -1362
rect -234 -1371 -230 -1344
rect -242 -1402 -238 -1391
rect -242 -1406 -230 -1402
rect -369 -1415 -346 -1410
rect -338 -1415 -294 -1410
rect -286 -1415 -242 -1410
rect -338 -1418 -334 -1415
rect -286 -1418 -282 -1415
rect -234 -1418 -230 -1406
rect -212 -1410 -207 -1344
rect -193 -1367 -190 -1362
rect -182 -1371 -178 -1344
rect -137 -1347 -133 -1344
rect -105 -1347 -101 -1344
rect -145 -1374 -141 -1367
rect -113 -1374 -109 -1367
rect -155 -1376 -91 -1374
rect -155 -1380 -153 -1376
rect -149 -1380 -129 -1376
rect -125 -1380 -121 -1376
rect -117 -1380 -97 -1376
rect -93 -1380 -91 -1376
rect -155 -1382 -91 -1380
rect -190 -1402 -186 -1391
rect -190 -1406 -178 -1402
rect -212 -1415 -190 -1410
rect -182 -1418 -178 -1406
rect -22 -1418 -17 -1313
rect 74 -1339 79 -1290
rect 111 -1308 115 -1307
rect 95 -1313 115 -1308
rect 119 -1312 123 -1307
rect 151 -1312 155 -1300
rect 189 -1312 193 -1300
rect 119 -1317 143 -1312
rect 151 -1317 181 -1312
rect 189 -1317 465 -1312
rect 119 -1319 123 -1317
rect 151 -1320 155 -1317
rect 189 -1320 193 -1317
rect 111 -1341 115 -1339
rect -9 -1379 0 -1376
rect -9 -1383 -6 -1379
rect -2 -1383 0 -1379
rect -9 -1386 0 -1383
rect -9 -1390 6 -1386
rect -9 -1401 0 -1390
rect 49 -1394 54 -1362
rect 74 -1368 79 -1344
rect 102 -1342 115 -1341
rect 102 -1346 103 -1342
rect 107 -1346 115 -1342
rect 102 -1347 115 -1346
rect 143 -1347 147 -1340
rect 181 -1347 185 -1340
rect 133 -1349 165 -1347
rect 133 -1353 135 -1349
rect 139 -1353 159 -1349
rect 163 -1353 165 -1349
rect 133 -1355 165 -1353
rect 171 -1349 203 -1347
rect 171 -1353 173 -1349
rect 177 -1353 197 -1349
rect 201 -1353 203 -1349
rect 171 -1355 203 -1353
rect 133 -1368 165 -1365
rect 58 -1373 111 -1368
rect 133 -1372 136 -1368
rect 140 -1372 158 -1368
rect 162 -1372 165 -1368
rect 58 -1386 63 -1373
rect 133 -1374 165 -1372
rect 342 -1368 412 -1365
rect 342 -1372 345 -1368
rect 349 -1372 405 -1368
rect 409 -1372 412 -1368
rect 342 -1374 412 -1372
rect 93 -1378 101 -1376
rect 93 -1382 95 -1378
rect 99 -1382 101 -1378
rect 143 -1380 147 -1374
rect 352 -1380 356 -1374
rect 390 -1380 394 -1374
rect 93 -1386 101 -1382
rect 86 -1390 101 -1386
rect 46 -1398 66 -1394
rect -9 -1405 -6 -1401
rect -2 -1405 0 -1401
rect -9 -1408 0 -1405
rect 58 -1409 63 -1398
rect 93 -1402 101 -1390
rect 93 -1406 95 -1402
rect 99 -1406 101 -1402
rect 111 -1403 115 -1401
rect 93 -1408 101 -1406
rect 104 -1407 115 -1403
rect 119 -1405 123 -1401
rect 58 -1414 83 -1409
rect 104 -1418 108 -1407
rect 119 -1410 132 -1405
rect 119 -1413 123 -1410
rect -79 -1423 108 -1418
rect -346 -1446 -342 -1438
rect -294 -1446 -290 -1438
rect -242 -1446 -238 -1438
rect -190 -1446 -186 -1438
rect -356 -1447 -168 -1446
rect -356 -1451 -329 -1447
rect -325 -1451 -277 -1447
rect -273 -1451 -225 -1447
rect -221 -1451 -173 -1447
rect -169 -1451 -168 -1447
rect -356 -1452 -168 -1451
rect -418 -1465 -356 -1460
rect -351 -1465 -304 -1460
rect -299 -1465 -250 -1460
rect -245 -1465 -198 -1460
rect -156 -1486 -92 -1483
rect -156 -1490 -153 -1486
rect -149 -1490 -131 -1486
rect -127 -1490 -121 -1486
rect -117 -1490 -99 -1486
rect -95 -1490 -92 -1486
rect -357 -1494 -169 -1491
rect -156 -1492 -92 -1490
rect -357 -1498 -354 -1494
rect -350 -1498 -332 -1494
rect -328 -1498 -302 -1494
rect -298 -1498 -280 -1494
rect -276 -1498 -250 -1494
rect -246 -1498 -228 -1494
rect -224 -1498 -198 -1494
rect -194 -1498 -176 -1494
rect -172 -1498 -169 -1494
rect -357 -1500 -169 -1498
rect -146 -1498 -142 -1492
rect -114 -1498 -110 -1492
rect -347 -1506 -343 -1500
rect -295 -1506 -291 -1500
rect -243 -1506 -239 -1500
rect -191 -1506 -187 -1500
rect -370 -1555 -347 -1550
rect -370 -1621 -365 -1555
rect -339 -1559 -335 -1546
rect -347 -1563 -335 -1559
rect -317 -1555 -295 -1550
rect -347 -1568 -343 -1563
rect -352 -1617 -347 -1612
rect -339 -1621 -335 -1608
rect -317 -1621 -312 -1555
rect -287 -1559 -283 -1546
rect -235 -1550 -231 -1546
rect -183 -1550 -179 -1546
rect -138 -1550 -134 -1538
rect -106 -1550 -102 -1538
rect -79 -1550 -74 -1423
rect -9 -1430 0 -1427
rect -9 -1434 -6 -1430
rect -2 -1434 0 -1430
rect -9 -1437 0 -1434
rect 58 -1437 63 -1423
rect 93 -1429 101 -1427
rect 93 -1433 95 -1429
rect 99 -1433 101 -1429
rect 93 -1437 101 -1433
rect -9 -1441 6 -1437
rect -9 -1452 0 -1441
rect 86 -1441 101 -1437
rect 46 -1449 66 -1445
rect -9 -1456 -6 -1452
rect -2 -1456 0 -1452
rect -9 -1459 0 -1456
rect 58 -1464 63 -1449
rect 93 -1453 101 -1441
rect 93 -1457 95 -1453
rect 99 -1457 101 -1453
rect 93 -1459 101 -1457
rect 127 -1432 132 -1410
rect 279 -1407 316 -1402
rect 151 -1432 155 -1420
rect 316 -1432 320 -1430
rect 111 -1464 115 -1433
rect 127 -1437 143 -1432
rect 151 -1437 283 -1432
rect 288 -1437 320 -1432
rect 460 -1400 465 -1317
rect 470 -1328 566 -1325
rect 470 -1332 499 -1328
rect 503 -1332 559 -1328
rect 563 -1332 566 -1328
rect 470 -1334 566 -1332
rect 470 -1370 474 -1334
rect 506 -1340 510 -1334
rect 544 -1340 548 -1334
rect 1332 -1353 1396 -1350
rect 1332 -1357 1335 -1353
rect 1339 -1357 1357 -1353
rect 1361 -1357 1367 -1353
rect 1371 -1357 1389 -1353
rect 1393 -1357 1396 -1353
rect 1131 -1361 1319 -1358
rect 1332 -1359 1396 -1357
rect 1131 -1365 1134 -1361
rect 1138 -1365 1156 -1361
rect 1160 -1365 1186 -1361
rect 1190 -1365 1208 -1361
rect 1212 -1365 1238 -1361
rect 1242 -1365 1260 -1361
rect 1264 -1365 1290 -1361
rect 1294 -1365 1312 -1361
rect 1316 -1365 1319 -1361
rect 1131 -1367 1319 -1365
rect 1342 -1365 1346 -1359
rect 1374 -1365 1378 -1359
rect 478 -1392 482 -1390
rect 514 -1392 518 -1380
rect 552 -1392 556 -1380
rect 1141 -1373 1145 -1367
rect 1193 -1373 1197 -1367
rect 1245 -1373 1249 -1367
rect 1297 -1373 1301 -1367
rect 478 -1397 506 -1392
rect 514 -1397 544 -1392
rect 552 -1397 809 -1392
rect 460 -1405 475 -1400
rect 478 -1405 482 -1397
rect 514 -1400 518 -1397
rect 552 -1400 556 -1397
rect 324 -1432 328 -1430
rect 360 -1432 364 -1420
rect 398 -1432 402 -1420
rect 324 -1437 352 -1432
rect 360 -1437 390 -1432
rect 398 -1437 470 -1432
rect 506 -1434 510 -1420
rect 544 -1434 548 -1420
rect 496 -1436 566 -1434
rect 151 -1440 155 -1437
rect 58 -1469 115 -1464
rect 324 -1445 328 -1437
rect 360 -1440 364 -1437
rect 398 -1440 402 -1437
rect 143 -1467 147 -1460
rect 496 -1440 498 -1436
rect 502 -1440 560 -1436
rect 564 -1440 566 -1436
rect 496 -1442 566 -1440
rect 133 -1469 165 -1467
rect 133 -1473 135 -1469
rect 139 -1473 159 -1469
rect 163 -1473 165 -1469
rect 133 -1475 165 -1473
rect 316 -1474 320 -1465
rect 352 -1474 356 -1460
rect 390 -1474 394 -1460
rect 306 -1476 412 -1474
rect 306 -1480 308 -1476
rect 312 -1480 406 -1476
rect 410 -1480 412 -1476
rect 306 -1482 412 -1480
rect 804 -1496 809 -1397
rect 1402 -1373 1434 -1370
rect 1402 -1377 1405 -1373
rect 1409 -1377 1427 -1373
rect 1431 -1377 1434 -1373
rect 1402 -1379 1434 -1377
rect 1412 -1385 1416 -1379
rect 819 -1424 915 -1421
rect 819 -1428 848 -1424
rect 852 -1428 908 -1424
rect 912 -1428 915 -1424
rect 819 -1430 915 -1428
rect 1118 -1422 1141 -1417
rect 819 -1466 823 -1430
rect 855 -1436 859 -1430
rect 893 -1436 897 -1430
rect 827 -1488 831 -1486
rect 863 -1488 867 -1476
rect 901 -1488 905 -1476
rect 1118 -1488 1123 -1422
rect 1149 -1426 1153 -1413
rect 1141 -1430 1153 -1426
rect 1171 -1422 1193 -1417
rect 1141 -1435 1145 -1430
rect 1136 -1484 1141 -1479
rect 1149 -1488 1153 -1475
rect 1171 -1488 1176 -1422
rect 1201 -1426 1205 -1413
rect 1253 -1417 1257 -1413
rect 1305 -1417 1309 -1413
rect 1350 -1417 1354 -1405
rect 1382 -1417 1386 -1405
rect 1420 -1417 1424 -1405
rect 1193 -1430 1205 -1426
rect 1223 -1422 1245 -1417
rect 1253 -1422 1297 -1417
rect 1305 -1422 1342 -1417
rect 1350 -1422 1374 -1417
rect 1382 -1422 1412 -1417
rect 1420 -1422 1434 -1417
rect 1193 -1435 1197 -1430
rect 1188 -1484 1193 -1479
rect 1201 -1488 1205 -1475
rect 1223 -1488 1228 -1422
rect 1242 -1445 1245 -1440
rect 1253 -1449 1257 -1422
rect 1245 -1480 1249 -1469
rect 1245 -1484 1257 -1480
rect 827 -1493 855 -1488
rect 863 -1493 893 -1488
rect 901 -1493 1141 -1488
rect 1149 -1493 1193 -1488
rect 1201 -1493 1245 -1488
rect 804 -1501 824 -1496
rect 827 -1501 831 -1493
rect 863 -1496 867 -1493
rect 901 -1496 905 -1493
rect 1149 -1496 1153 -1493
rect 1201 -1496 1205 -1493
rect 1253 -1496 1257 -1484
rect 1275 -1488 1280 -1422
rect 1294 -1445 1297 -1440
rect 1305 -1449 1309 -1422
rect 1350 -1425 1354 -1422
rect 1382 -1425 1386 -1422
rect 1420 -1425 1424 -1422
rect 1412 -1442 1416 -1435
rect 1402 -1444 1434 -1442
rect 1342 -1452 1346 -1445
rect 1374 -1452 1378 -1445
rect 1402 -1448 1404 -1444
rect 1408 -1448 1428 -1444
rect 1432 -1448 1434 -1444
rect 1402 -1450 1434 -1448
rect 1332 -1454 1396 -1452
rect 1332 -1458 1334 -1454
rect 1338 -1458 1358 -1454
rect 1362 -1458 1366 -1454
rect 1370 -1458 1390 -1454
rect 1394 -1458 1396 -1454
rect 1332 -1460 1396 -1458
rect 1297 -1480 1301 -1469
rect 1297 -1484 1309 -1480
rect 1275 -1493 1297 -1488
rect 1305 -1496 1309 -1484
rect 342 -1512 412 -1509
rect 342 -1516 345 -1512
rect 349 -1516 405 -1512
rect 409 -1516 412 -1512
rect 342 -1518 412 -1516
rect 352 -1524 356 -1518
rect 390 -1524 394 -1518
rect -295 -1563 -283 -1559
rect -265 -1555 -243 -1550
rect -235 -1555 -191 -1550
rect -183 -1555 -146 -1550
rect -138 -1555 -114 -1550
rect -106 -1555 -74 -1550
rect 288 -1551 316 -1546
rect -295 -1568 -291 -1563
rect -300 -1617 -295 -1612
rect -287 -1621 -283 -1608
rect -265 -1621 -260 -1555
rect -246 -1578 -243 -1573
rect -235 -1582 -231 -1555
rect -243 -1613 -239 -1602
rect -243 -1617 -231 -1613
rect -370 -1626 -347 -1621
rect -339 -1626 -295 -1621
rect -287 -1626 -243 -1621
rect -339 -1629 -335 -1626
rect -287 -1629 -283 -1626
rect -235 -1629 -231 -1617
rect -213 -1621 -208 -1555
rect -194 -1578 -191 -1573
rect -183 -1582 -179 -1555
rect -138 -1558 -134 -1555
rect -106 -1558 -102 -1555
rect 316 -1576 320 -1574
rect -146 -1585 -142 -1578
rect -114 -1585 -110 -1578
rect 270 -1581 320 -1576
rect 809 -1533 819 -1528
rect 855 -1530 859 -1516
rect 893 -1530 897 -1516
rect 1141 -1524 1145 -1516
rect 1193 -1524 1197 -1516
rect 1245 -1524 1249 -1516
rect 1297 -1524 1301 -1516
rect 1131 -1525 1319 -1524
rect 1131 -1529 1158 -1525
rect 1162 -1529 1210 -1525
rect 1214 -1529 1262 -1525
rect 1266 -1529 1314 -1525
rect 1318 -1529 1319 -1525
rect 1131 -1530 1319 -1529
rect 845 -1532 915 -1530
rect 471 -1542 541 -1539
rect 471 -1546 474 -1542
rect 478 -1546 534 -1542
rect 538 -1546 541 -1542
rect 471 -1548 541 -1546
rect 324 -1576 328 -1574
rect 360 -1576 364 -1564
rect 398 -1576 402 -1564
rect 481 -1554 485 -1548
rect 519 -1554 523 -1548
rect 324 -1581 352 -1576
rect 360 -1581 390 -1576
rect 398 -1581 445 -1576
rect -156 -1587 -92 -1585
rect -156 -1591 -154 -1587
rect -150 -1591 -130 -1587
rect -126 -1591 -122 -1587
rect -118 -1591 -98 -1587
rect -94 -1591 -92 -1587
rect 324 -1589 328 -1581
rect 360 -1584 364 -1581
rect 398 -1584 402 -1581
rect -156 -1593 -92 -1591
rect -191 -1613 -187 -1602
rect -191 -1617 -179 -1613
rect -213 -1626 -191 -1621
rect -183 -1629 -179 -1617
rect 316 -1618 320 -1609
rect 352 -1618 356 -1604
rect 390 -1618 394 -1604
rect 445 -1606 449 -1604
rect 425 -1611 449 -1606
rect 453 -1606 457 -1604
rect 489 -1606 493 -1594
rect 527 -1606 531 -1594
rect 579 -1603 675 -1600
rect 453 -1611 481 -1606
rect 489 -1611 519 -1606
rect 527 -1611 574 -1606
rect 306 -1620 412 -1618
rect 306 -1624 308 -1620
rect 312 -1624 406 -1620
rect 410 -1624 412 -1620
rect 306 -1626 412 -1624
rect 425 -1641 431 -1611
rect 453 -1619 457 -1611
rect 489 -1614 493 -1611
rect 527 -1614 531 -1611
rect 261 -1646 431 -1641
rect 445 -1648 449 -1639
rect 481 -1648 485 -1634
rect 519 -1648 523 -1634
rect -347 -1657 -343 -1649
rect -295 -1657 -291 -1649
rect -243 -1657 -239 -1649
rect -191 -1657 -187 -1649
rect 435 -1650 541 -1648
rect 435 -1654 437 -1650
rect 441 -1654 535 -1650
rect 539 -1654 541 -1650
rect 435 -1656 541 -1654
rect -357 -1658 -169 -1657
rect -357 -1662 -330 -1658
rect -326 -1662 -278 -1658
rect -274 -1662 -226 -1658
rect -222 -1662 -174 -1658
rect -170 -1662 -169 -1658
rect -357 -1663 -169 -1662
rect -418 -1676 -357 -1671
rect -352 -1676 -305 -1671
rect -300 -1676 -251 -1671
rect -246 -1676 -199 -1671
rect 569 -1675 574 -1611
rect 579 -1607 608 -1603
rect 612 -1607 668 -1603
rect 672 -1607 675 -1603
rect 579 -1609 675 -1607
rect 579 -1645 583 -1609
rect 615 -1615 619 -1609
rect 653 -1615 657 -1609
rect 587 -1667 591 -1665
rect 623 -1667 627 -1655
rect 661 -1667 665 -1655
rect 587 -1672 615 -1667
rect 623 -1672 653 -1667
rect 661 -1672 698 -1667
rect 345 -1682 415 -1679
rect 569 -1680 584 -1675
rect 587 -1680 591 -1672
rect 623 -1675 627 -1672
rect 661 -1675 665 -1672
rect 345 -1686 348 -1682
rect 352 -1686 408 -1682
rect 412 -1686 415 -1682
rect 345 -1688 415 -1686
rect 355 -1694 359 -1688
rect 393 -1694 397 -1688
rect 288 -1721 319 -1716
rect 319 -1746 323 -1744
rect 270 -1751 323 -1746
rect 476 -1712 546 -1709
rect 476 -1716 479 -1712
rect 483 -1716 539 -1712
rect 543 -1716 546 -1712
rect 476 -1718 546 -1716
rect 569 -1712 579 -1707
rect 615 -1709 619 -1695
rect 653 -1709 657 -1695
rect 605 -1711 675 -1709
rect 327 -1746 331 -1744
rect 363 -1746 367 -1734
rect 401 -1746 405 -1734
rect 486 -1724 490 -1718
rect 524 -1724 528 -1718
rect 327 -1751 355 -1746
rect 363 -1751 393 -1746
rect 401 -1751 450 -1746
rect 327 -1759 331 -1751
rect 363 -1754 367 -1751
rect 401 -1754 405 -1751
rect 319 -1788 323 -1779
rect 355 -1788 359 -1774
rect 393 -1788 397 -1774
rect 450 -1776 454 -1774
rect 420 -1781 454 -1776
rect 458 -1776 462 -1774
rect 494 -1776 498 -1764
rect 532 -1776 536 -1764
rect 569 -1776 574 -1712
rect 605 -1715 607 -1711
rect 611 -1715 669 -1711
rect 673 -1715 675 -1711
rect 605 -1717 675 -1715
rect 458 -1781 486 -1776
rect 494 -1781 524 -1776
rect 532 -1781 574 -1776
rect 309 -1790 415 -1788
rect 309 -1794 311 -1790
rect 315 -1794 409 -1790
rect 413 -1794 415 -1790
rect 309 -1796 415 -1794
rect 345 -1826 415 -1823
rect 345 -1830 348 -1826
rect 352 -1830 408 -1826
rect 412 -1830 415 -1826
rect 345 -1832 415 -1830
rect 355 -1838 359 -1832
rect 393 -1838 397 -1832
rect 252 -1865 319 -1860
rect 319 -1890 323 -1888
rect 243 -1895 323 -1890
rect 327 -1890 331 -1888
rect 363 -1890 367 -1878
rect 401 -1890 405 -1878
rect 420 -1890 425 -1781
rect 458 -1789 462 -1781
rect 494 -1784 498 -1781
rect 532 -1784 536 -1781
rect 450 -1818 454 -1809
rect 486 -1818 490 -1804
rect 524 -1818 528 -1804
rect 440 -1820 546 -1818
rect 440 -1824 442 -1820
rect 446 -1824 540 -1820
rect 544 -1824 546 -1820
rect 440 -1826 546 -1824
rect 693 -1864 698 -1672
rect 708 -1792 804 -1789
rect 708 -1796 737 -1792
rect 741 -1796 797 -1792
rect 801 -1796 804 -1792
rect 708 -1798 804 -1796
rect 708 -1834 712 -1798
rect 744 -1804 748 -1798
rect 782 -1804 786 -1798
rect 716 -1856 720 -1854
rect 752 -1856 756 -1844
rect 790 -1856 794 -1844
rect 809 -1856 814 -1533
rect 845 -1536 847 -1532
rect 851 -1536 909 -1532
rect 913 -1536 915 -1532
rect 845 -1538 915 -1536
rect 1105 -1543 1131 -1538
rect 1136 -1543 1183 -1538
rect 1188 -1543 1237 -1538
rect 1242 -1543 1289 -1538
rect 716 -1861 744 -1856
rect 752 -1861 782 -1856
rect 790 -1861 814 -1856
rect 693 -1869 713 -1864
rect 716 -1869 720 -1861
rect 752 -1864 756 -1861
rect 790 -1864 794 -1861
rect 327 -1895 355 -1890
rect 363 -1895 393 -1890
rect 401 -1895 425 -1890
rect 327 -1903 331 -1895
rect 363 -1898 367 -1895
rect 401 -1898 405 -1895
rect 693 -1901 708 -1896
rect 744 -1898 748 -1884
rect 782 -1898 786 -1884
rect 734 -1900 804 -1898
rect 319 -1932 323 -1923
rect 355 -1932 359 -1918
rect 393 -1932 397 -1918
rect 309 -1934 415 -1932
rect 309 -1938 311 -1934
rect 315 -1938 409 -1934
rect 413 -1938 415 -1934
rect 309 -1940 415 -1938
rect 345 -1953 415 -1950
rect 345 -1957 348 -1953
rect 352 -1957 408 -1953
rect 412 -1957 415 -1953
rect 345 -1959 415 -1957
rect 355 -1965 359 -1959
rect 393 -1965 397 -1959
rect 288 -1992 319 -1987
rect 319 -2017 323 -2015
rect 270 -2022 323 -2017
rect 476 -1983 546 -1980
rect 476 -1987 479 -1983
rect 483 -1987 539 -1983
rect 543 -1987 546 -1983
rect 476 -1989 546 -1987
rect 327 -2017 331 -2015
rect 363 -2017 367 -2005
rect 401 -2017 405 -2005
rect 486 -1995 490 -1989
rect 524 -1995 528 -1989
rect 327 -2022 355 -2017
rect 363 -2022 393 -2017
rect 401 -2022 450 -2017
rect 327 -2030 331 -2022
rect 363 -2025 367 -2022
rect 401 -2025 405 -2022
rect 319 -2059 323 -2050
rect 355 -2059 359 -2045
rect 393 -2059 397 -2045
rect 450 -2047 454 -2045
rect 420 -2052 454 -2047
rect 611 -2013 681 -2010
rect 611 -2017 614 -2013
rect 618 -2017 674 -2013
rect 678 -2017 681 -2013
rect 611 -2019 681 -2017
rect 458 -2047 462 -2045
rect 494 -2047 498 -2035
rect 532 -2047 536 -2035
rect 621 -2025 625 -2019
rect 659 -2025 663 -2019
rect 458 -2052 486 -2047
rect 494 -2052 524 -2047
rect 532 -2052 585 -2047
rect 309 -2061 415 -2059
rect 309 -2065 311 -2061
rect 315 -2065 409 -2061
rect 413 -2065 415 -2061
rect 309 -2067 415 -2065
rect 345 -2097 415 -2094
rect 345 -2101 348 -2097
rect 352 -2101 408 -2097
rect 412 -2101 415 -2097
rect 345 -2103 415 -2101
rect 355 -2109 359 -2103
rect 393 -2109 397 -2103
rect 252 -2136 319 -2131
rect 319 -2161 323 -2159
rect 234 -2166 323 -2161
rect 327 -2161 331 -2159
rect 363 -2161 367 -2149
rect 401 -2161 405 -2149
rect 420 -2161 425 -2052
rect 458 -2060 462 -2052
rect 494 -2055 498 -2052
rect 532 -2055 536 -2052
rect 450 -2089 454 -2080
rect 486 -2089 490 -2075
rect 524 -2089 528 -2075
rect 585 -2077 589 -2075
rect 558 -2082 589 -2077
rect 593 -2077 597 -2075
rect 629 -2077 633 -2065
rect 667 -2077 671 -2065
rect 693 -2077 698 -1901
rect 734 -1904 736 -1900
rect 740 -1904 798 -1900
rect 802 -1904 804 -1900
rect 734 -1906 804 -1904
rect 593 -2082 621 -2077
rect 629 -2082 659 -2077
rect 667 -2082 698 -2077
rect 440 -2091 546 -2089
rect 440 -2095 442 -2091
rect 446 -2095 540 -2091
rect 544 -2095 546 -2091
rect 440 -2097 546 -2095
rect 327 -2166 355 -2161
rect 363 -2166 393 -2161
rect 401 -2166 425 -2161
rect 327 -2174 331 -2166
rect 363 -2169 367 -2166
rect 401 -2169 405 -2166
rect 319 -2203 323 -2194
rect 355 -2203 359 -2189
rect 393 -2203 397 -2189
rect 309 -2205 415 -2203
rect 309 -2209 311 -2205
rect 315 -2209 409 -2205
rect 413 -2209 415 -2205
rect 309 -2211 415 -2209
rect 558 -2220 563 -2082
rect 593 -2090 597 -2082
rect 629 -2085 633 -2082
rect 667 -2085 671 -2082
rect 585 -2119 589 -2110
rect 621 -2119 625 -2105
rect 659 -2119 663 -2105
rect 575 -2121 681 -2119
rect 575 -2125 577 -2121
rect 581 -2125 675 -2121
rect 679 -2125 681 -2121
rect 575 -2127 681 -2125
rect 225 -2225 563 -2220
<< m2contact >>
rect -423 363 -418 368
rect 1100 363 1105 368
rect 220 280 225 285
rect 229 230 234 235
rect -354 117 -349 122
rect 1132 225 1137 230
rect 1184 225 1189 230
rect 1238 264 1243 269
rect 1290 264 1295 269
rect -302 117 -297 122
rect -248 156 -243 161
rect -196 156 -191 161
rect 1100 166 1105 171
rect 1132 166 1137 171
rect 1184 166 1189 171
rect 1238 166 1243 171
rect 1290 166 1295 171
rect -80 69 -75 74
rect 58 95 63 100
rect -423 58 -418 63
rect -354 58 -349 63
rect -302 58 -297 63
rect -248 58 -243 63
rect -196 58 -191 63
rect 90 95 95 100
rect 238 91 243 96
rect 74 69 79 74
rect -355 -94 -350 -89
rect -303 -94 -298 -89
rect -249 -55 -244 -50
rect -197 -55 -192 -50
rect 229 1 234 6
rect 220 -29 225 -24
rect 889 49 894 54
rect 1131 25 1136 30
rect 1183 25 1188 30
rect 1237 64 1242 69
rect 1289 64 1294 69
rect 1100 -34 1105 -29
rect 1131 -34 1136 -29
rect 1183 -34 1188 -29
rect 1237 -34 1242 -29
rect 1289 -34 1294 -29
rect 247 -86 252 -81
rect 464 -86 469 -81
rect -423 -153 -418 -148
rect -355 -153 -350 -148
rect -303 -153 -298 -148
rect -249 -153 -244 -148
rect -197 -153 -192 -148
rect -363 -298 -358 -293
rect 58 -195 63 -190
rect -99 -236 -94 -231
rect -311 -298 -306 -293
rect -257 -259 -252 -254
rect -205 -259 -200 -254
rect 90 -195 95 -190
rect 256 -199 261 -194
rect 74 -236 79 -231
rect -423 -357 -418 -352
rect -363 -357 -358 -352
rect -311 -357 -306 -352
rect -257 -357 -252 -352
rect -205 -357 -200 -352
rect -364 -509 -359 -504
rect 238 -289 243 -284
rect 247 -319 252 -314
rect 220 -415 225 -410
rect 229 -445 234 -440
rect -312 -509 -307 -504
rect -258 -470 -253 -465
rect -206 -470 -201 -465
rect 889 -363 894 -358
rect 1130 -374 1135 -369
rect 1182 -374 1187 -369
rect 1236 -335 1241 -330
rect 1288 -335 1293 -330
rect 1100 -433 1105 -428
rect 1130 -433 1135 -428
rect 1182 -433 1187 -428
rect 1236 -433 1241 -428
rect 1288 -433 1293 -428
rect 247 -511 252 -505
rect 265 -533 270 -528
rect 645 -533 650 -528
rect -423 -568 -418 -563
rect -364 -568 -359 -563
rect -312 -568 -307 -563
rect -258 -568 -253 -563
rect -206 -568 -201 -563
rect -369 -704 -364 -699
rect 58 -612 63 -607
rect -103 -642 -98 -637
rect -317 -704 -312 -699
rect -263 -665 -258 -660
rect -211 -665 -206 -660
rect 90 -612 95 -607
rect 274 -616 279 -611
rect 74 -642 79 -637
rect -423 -763 -418 -758
rect -369 -763 -364 -758
rect -317 -763 -312 -758
rect -263 -763 -258 -758
rect -211 -763 -206 -758
rect -370 -915 -365 -910
rect 256 -706 261 -701
rect 265 -736 270 -731
rect 238 -850 243 -845
rect -318 -915 -313 -910
rect -264 -876 -259 -871
rect -212 -876 -207 -871
rect 247 -880 252 -875
rect 265 -945 270 -940
rect 890 -795 895 -790
rect 1130 -788 1135 -783
rect 1182 -788 1187 -783
rect 1236 -749 1241 -744
rect 1288 -749 1293 -744
rect 1100 -847 1105 -842
rect 1130 -847 1135 -842
rect 1182 -847 1187 -842
rect 1236 -847 1241 -842
rect 1288 -847 1293 -842
rect -423 -974 -418 -969
rect -370 -974 -365 -969
rect -318 -974 -313 -969
rect -264 -974 -259 -969
rect -212 -974 -207 -969
rect 220 -1020 225 -1015
rect 229 -1050 234 -1045
rect 247 -1164 252 -1159
rect 265 -1194 270 -1189
rect 283 -1249 288 -1244
rect 853 -1249 858 -1244
rect -356 -1406 -351 -1401
rect 58 -1313 63 -1308
rect -93 -1344 -88 -1339
rect -304 -1406 -299 -1401
rect -250 -1367 -245 -1362
rect -198 -1367 -193 -1362
rect 90 -1313 95 -1308
rect 74 -1344 79 -1339
rect -423 -1465 -418 -1460
rect -356 -1465 -351 -1460
rect -304 -1465 -299 -1460
rect -250 -1465 -245 -1460
rect -198 -1465 -193 -1460
rect -357 -1617 -352 -1612
rect 274 -1407 279 -1402
rect 283 -1437 288 -1432
rect 1131 -1484 1136 -1479
rect 1183 -1484 1188 -1479
rect 1237 -1445 1242 -1440
rect 1289 -1445 1294 -1440
rect 283 -1551 288 -1546
rect -305 -1617 -300 -1612
rect -251 -1578 -246 -1573
rect -199 -1578 -194 -1573
rect 265 -1581 270 -1576
rect 256 -1646 261 -1641
rect -423 -1676 -418 -1671
rect -357 -1676 -352 -1671
rect -305 -1676 -300 -1671
rect -251 -1676 -246 -1671
rect -199 -1676 -194 -1671
rect 283 -1721 288 -1716
rect 265 -1751 270 -1746
rect 247 -1865 252 -1860
rect 238 -1895 243 -1890
rect 1100 -1543 1105 -1538
rect 1131 -1543 1136 -1538
rect 1183 -1543 1188 -1538
rect 1237 -1543 1242 -1538
rect 1289 -1543 1294 -1538
rect 283 -1992 288 -1987
rect 265 -2022 270 -2017
rect 247 -2136 252 -2131
rect 229 -2166 234 -2161
rect 220 -2225 225 -2220
<< metal2 >>
rect -423 63 -418 363
rect -354 63 -349 117
rect -302 63 -297 117
rect -248 63 -243 156
rect -196 63 -191 156
rect 63 95 90 100
rect -75 69 74 74
rect -423 -148 -418 58
rect 220 -24 225 280
rect -355 -148 -350 -94
rect -303 -148 -298 -94
rect -249 -148 -244 -55
rect -197 -148 -192 -55
rect -423 -352 -418 -153
rect 63 -195 90 -190
rect -94 -236 74 -231
rect -363 -352 -358 -298
rect -311 -352 -306 -298
rect -257 -352 -252 -259
rect -205 -352 -200 -259
rect -423 -563 -418 -357
rect 220 -410 225 -29
rect -364 -563 -359 -509
rect -312 -563 -307 -509
rect -258 -563 -253 -470
rect -206 -563 -201 -470
rect -423 -758 -418 -568
rect 63 -612 90 -607
rect -98 -642 74 -637
rect -369 -758 -364 -704
rect -317 -758 -312 -704
rect -263 -758 -258 -665
rect -211 -758 -206 -665
rect -423 -969 -418 -763
rect -370 -969 -365 -915
rect -318 -969 -313 -915
rect -264 -969 -259 -876
rect -212 -969 -207 -876
rect -423 -1460 -418 -974
rect 220 -1015 225 -415
rect 63 -1313 90 -1308
rect -88 -1344 74 -1339
rect -356 -1460 -351 -1406
rect -304 -1460 -299 -1406
rect -250 -1460 -245 -1367
rect -198 -1460 -193 -1367
rect -423 -1671 -418 -1465
rect -357 -1671 -352 -1617
rect -305 -1671 -300 -1617
rect -251 -1671 -246 -1578
rect -199 -1671 -194 -1578
rect 220 -2220 225 -1020
rect 229 6 234 230
rect 1100 171 1105 363
rect 1132 171 1137 225
rect 1184 171 1189 225
rect 1238 171 1243 264
rect 1290 171 1295 264
rect 229 -440 234 1
rect 229 -1045 234 -445
rect 229 -2161 234 -1050
rect 238 -284 243 91
rect 464 49 889 54
rect 464 -81 469 49
rect 238 -845 243 -289
rect 238 -1890 243 -850
rect 1100 -29 1105 166
rect 1131 -29 1136 25
rect 1183 -29 1188 25
rect 1237 -29 1242 64
rect 1289 -29 1294 64
rect 247 -314 252 -86
rect 247 -505 252 -319
rect 247 -875 252 -511
rect 247 -1159 252 -880
rect 247 -1860 252 -1164
rect 256 -701 261 -199
rect 645 -363 889 -358
rect 645 -528 650 -363
rect 256 -1641 261 -706
rect 1100 -428 1105 -34
rect 1130 -428 1135 -374
rect 1182 -428 1187 -374
rect 1236 -428 1241 -335
rect 1288 -428 1293 -335
rect 265 -731 270 -533
rect 265 -940 270 -736
rect 265 -1189 270 -945
rect 265 -1576 270 -1194
rect 274 -1402 279 -616
rect 853 -795 890 -790
rect 853 -1244 858 -795
rect 1100 -842 1105 -433
rect 1130 -842 1135 -788
rect 1182 -842 1187 -788
rect 1236 -842 1241 -749
rect 1288 -842 1293 -749
rect 247 -2131 252 -1865
rect 265 -1746 270 -1581
rect 265 -2017 270 -1751
rect 283 -1432 288 -1249
rect 283 -1546 288 -1437
rect 1100 -1538 1105 -847
rect 1131 -1538 1136 -1484
rect 1183 -1538 1188 -1484
rect 1237 -1538 1242 -1445
rect 1289 -1538 1294 -1445
rect 283 -1716 288 -1551
rect 283 -1987 288 -1721
<< labels >>
rlabel metal1 -5 -35 -5 -35 3 vdd
rlabel metal1 97 -34 97 -34 7 gnd
rlabel metal1 97 17 97 17 7 gnd
rlabel metal1 -5 16 -5 16 3 vdd
rlabel metal1 149 39 149 39 5 vdd
rlabel metal1 149 159 149 159 5 vdd
rlabel metal1 148 57 148 57 1 gnd
rlabel metal1 187 159 187 159 5 vdd
rlabel metal1 186 57 186 57 1 gnd
rlabel metal1 111 64 111 64 1 gnd
rlabel metal1 148 -63 148 -63 1 gnd
rlabel metal1 60 0 60 0 1 a0_not
rlabel metal1 85 -59 85 -59 1 b0_not
rlabel metal1 130 -13 130 -13 1 p0_not
rlabel metal1 160 -26 160 -26 1 p0
rlabel metal1 135 94 135 94 1 g0_mid
rlabel metal1 169 94 169 94 1 g0_not
rlabel metal1 200 94 200 94 1 g0
rlabel metal1 -5 -325 -5 -325 3 vdd
rlabel metal1 97 -324 97 -324 7 gnd
rlabel metal1 97 -273 97 -273 7 gnd
rlabel metal1 -5 -274 -5 -274 3 vdd
rlabel metal1 149 -251 149 -251 5 vdd
rlabel metal1 148 -353 148 -353 1 gnd
rlabel metal1 149 -131 149 -131 5 vdd
rlabel metal1 148 -233 148 -233 1 gnd
rlabel metal1 187 -131 187 -131 5 vdd
rlabel metal1 186 -233 186 -233 1 gnd
rlabel metal1 111 -226 111 -226 1 gnd
rlabel metal1 200 -196 200 -196 1 g1
rlabel metal1 169 -196 169 -196 1 g1_not
rlabel metal1 135 -196 135 -196 1 g1_mid
rlabel metal1 60 -290 60 -290 1 a1_not
rlabel metal1 85 -349 85 -349 1 b1_not
rlabel metal1 130 -303 130 -303 1 p1_not
rlabel metal1 160 -316 160 -316 1 p1
rlabel metal1 111 -643 111 -643 1 gnd
rlabel metal1 186 -650 186 -650 1 gnd
rlabel metal1 187 -548 187 -548 5 vdd
rlabel metal1 148 -650 148 -650 1 gnd
rlabel metal1 149 -548 149 -548 5 vdd
rlabel metal1 148 -770 148 -770 1 gnd
rlabel metal1 149 -668 149 -668 5 vdd
rlabel metal1 -5 -691 -5 -691 3 vdd
rlabel metal1 97 -690 97 -690 7 gnd
rlabel metal1 97 -741 97 -741 7 gnd
rlabel metal1 -5 -742 -5 -742 3 vdd
rlabel metal1 135 -613 135 -613 1 g2_mid
rlabel metal1 169 -613 169 -613 1 g2_not
rlabel metal1 200 -613 200 -613 1 g2
rlabel metal1 160 -733 160 -733 1 p2
rlabel metal1 130 -720 130 -720 1 p2_not
rlabel metal1 60 -707 60 -707 1 a2_not
rlabel metal1 85 -766 85 -766 1 b2_not
rlabel metal1 365 -27 365 -27 1 w1
rlabel metal1 333 38 333 38 5 vdd
rlabel metal1 318 -70 318 -70 1 gnd
rlabel metal1 424 58 424 58 1 gnd
rlabel metal1 439 166 439 166 5 vdd
rlabel metal1 473 101 473 101 1 c1
rlabel metal1 413 -252 413 -252 5 vdd
rlabel metal1 398 -360 398 -360 1 gnd
rlabel metal1 255 -27 255 -27 1 p0
rlabel metal1 249 3 249 3 1 c0
rlabel metal1 328 -286 328 -286 1 g0
rlabel metal1 328 -317 328 -317 1 p1
rlabel metal1 326 -486 326 -486 1 gnd
rlabel metal1 341 -378 341 -378 5 vdd
rlabel metal1 270 -413 270 -413 1 p0
rlabel metal1 270 -443 270 -443 1 c0
rlabel metal1 455 -516 455 -516 1 gnd
rlabel metal1 470 -408 470 -408 5 vdd
rlabel metal1 513 -473 513 -473 1 p1p0c0
rlabel metal1 457 -256 457 -256 1 p1g0
rlabel metal1 501 -232 501 -232 1 gnd
rlabel metal1 516 -124 516 -124 5 vdd
rlabel metal1 365 -669 365 -669 5 vdd
rlabel metal1 350 -777 350 -777 1 gnd
rlabel metal1 350 -921 350 -921 1 gnd
rlabel metal1 365 -813 365 -813 5 vdd
rlabel metal1 479 -951 479 -951 1 gnd
rlabel metal1 494 -843 494 -843 5 vdd
rlabel metal1 368 -983 368 -983 5 vdd
rlabel metal1 353 -1091 353 -1091 1 gnd
rlabel metal1 368 -1127 368 -1127 5 vdd
rlabel metal1 353 -1235 353 -1235 1 gnd
rlabel nwell 187 -1306 187 -1306 5 vdd
rlabel nwell 149 -1306 149 -1306 5 vdd
rlabel metal1 484 -1121 484 -1121 1 gnd
rlabel metal1 499 -1013 499 -1013 5 vdd
rlabel metal1 673 -541 673 -541 5 vdd
rlabel metal1 658 -649 658 -649 1 gnd
rlabel metal1 669 -897 669 -897 5 vdd
rlabel metal1 654 -1005 654 -1005 1 gnd
rlabel metal1 840 -678 840 -678 5 vdd
rlabel metal1 825 -786 825 -786 1 gnd
rlabel metal1 667 -310 667 -310 1 c2
rlabel metal1 621 -354 621 -354 1 gnd
rlabel metal1 636 -246 636 -246 5 vdd
rlabel metal1 873 -743 873 -743 7 c3
rlabel metal1 111 -1344 111 -1344 1 gnd
rlabel metal1 186 -1351 186 -1351 1 gnd
rlabel metal1 148 -1351 148 -1351 1 gnd
rlabel metal1 148 -1471 148 -1471 1 gnd
rlabel metal1 149 -1369 149 -1369 5 vdd
rlabel metal1 -5 -1392 -5 -1392 3 vdd
rlabel metal1 97 -1391 97 -1391 7 gnd
rlabel metal1 97 -1442 97 -1442 7 gnd
rlabel metal1 -5 -1443 -5 -1443 3 vdd
rlabel metal1 135 -1314 135 -1314 1 g3_mid
rlabel metal1 169 -1314 169 -1314 1 g3_not
rlabel metal1 200 -1314 200 -1314 1 g3
rlabel metal1 160 -1434 160 -1434 1 p3
rlabel metal1 60 -1408 60 -1408 1 a3_not
rlabel metal1 85 -1467 85 -1467 1 b3_not
rlabel metal1 130 -1421 130 -1421 1 p3_not
rlabel metal1 149 -1249 149 -1249 5 vdd
rlabel metal1 187 -1249 187 -1249 5 vdd
rlabel metal1 511 -1714 511 -1714 5 vdd
rlabel metal1 496 -1822 496 -1822 1 gnd
rlabel metal1 365 -1936 365 -1936 1 gnd
rlabel metal1 380 -1828 380 -1828 5 vdd
rlabel metal1 365 -1792 365 -1792 1 gnd
rlabel metal1 380 -1684 380 -1684 5 vdd
rlabel metal1 506 -1544 506 -1544 5 vdd
rlabel metal1 491 -1652 491 -1652 1 gnd
rlabel metal1 377 -1514 377 -1514 5 vdd
rlabel metal1 362 -1622 362 -1622 1 gnd
rlabel metal1 362 -1478 362 -1478 1 gnd
rlabel metal1 377 -1370 377 -1370 5 vdd
rlabel metal1 511 -1985 511 -1985 5 vdd
rlabel metal1 496 -2093 496 -2093 1 gnd
rlabel metal1 365 -2207 365 -2207 1 gnd
rlabel metal1 380 -2099 380 -2099 5 vdd
rlabel metal1 365 -2063 365 -2063 1 gnd
rlabel metal1 380 -1955 380 -1955 5 vdd
rlabel metal1 646 -2015 646 -2015 5 vdd
rlabel metal1 631 -2123 631 -2123 1 gnd
rlabel metal1 516 -1438 516 -1438 1 gnd
rlabel metal1 531 -1330 531 -1330 5 vdd
rlabel metal1 640 -1605 640 -1605 5 vdd
rlabel metal1 625 -1713 625 -1713 1 gnd
rlabel metal1 769 -1794 769 -1794 5 vdd
rlabel metal1 754 -1902 754 -1902 1 gnd
rlabel metal1 865 -1534 865 -1534 1 gnd
rlabel metal1 880 -1426 880 -1426 5 vdd
rlabel metal1 -338 239 -338 239 5 vdd
rlabel metal1 -338 74 -338 74 1 gnd
rlabel metal1 -286 239 -286 239 5 vdd
rlabel metal1 -286 74 -286 74 1 gnd
rlabel metal1 -234 74 -234 74 1 gnd
rlabel metal1 -234 239 -234 239 5 vdd
rlabel metal1 -182 74 -182 74 1 gnd
rlabel metal1 -182 239 -182 239 5 vdd
rlabel metal1 -106 145 -106 145 1 gnd
rlabel metal1 -105 247 -105 247 5 vdd
rlabel metal1 -138 145 -138 145 1 gnd
rlabel metal1 -137 247 -137 247 5 vdd
rlabel metal1 -339 28 -339 28 5 vdd
rlabel metal1 -339 -137 -339 -137 1 gnd
rlabel metal1 -287 28 -287 28 5 vdd
rlabel metal1 -287 -137 -287 -137 1 gnd
rlabel metal1 -235 -137 -235 -137 1 gnd
rlabel metal1 -235 28 -235 28 5 vdd
rlabel metal1 -183 -137 -183 -137 1 gnd
rlabel metal1 -183 28 -183 28 5 vdd
rlabel metal1 -107 -66 -107 -66 1 gnd
rlabel metal1 -106 36 -106 36 5 vdd
rlabel metal1 -139 -66 -139 -66 1 gnd
rlabel metal1 -138 36 -138 36 5 vdd
rlabel metal1 -365 151 -365 151 3 a0
rlabel metal1 -365 -61 -365 -61 3 b0
rlabel metal1 -77 128 -77 128 1 a0mid
rlabel metal1 -67 -30 -67 -30 1 b0mid
rlabel metal1 -347 -176 -347 -176 5 vdd
rlabel metal1 -347 -341 -347 -341 1 gnd
rlabel metal1 -295 -176 -295 -176 5 vdd
rlabel metal1 -295 -341 -295 -341 1 gnd
rlabel metal1 -243 -341 -243 -341 1 gnd
rlabel metal1 -243 -176 -243 -176 5 vdd
rlabel metal1 -191 -341 -191 -341 1 gnd
rlabel metal1 -191 -176 -191 -176 5 vdd
rlabel metal1 -115 -270 -115 -270 1 gnd
rlabel metal1 -114 -168 -114 -168 5 vdd
rlabel metal1 -147 -270 -147 -270 1 gnd
rlabel metal1 -146 -168 -146 -168 5 vdd
rlabel metal1 -348 -387 -348 -387 5 vdd
rlabel metal1 -348 -552 -348 -552 1 gnd
rlabel metal1 -296 -387 -296 -387 5 vdd
rlabel metal1 -296 -552 -296 -552 1 gnd
rlabel metal1 -244 -552 -244 -552 1 gnd
rlabel metal1 -244 -387 -244 -387 5 vdd
rlabel metal1 -192 -552 -192 -552 1 gnd
rlabel metal1 -192 -387 -192 -387 5 vdd
rlabel metal1 -116 -481 -116 -481 1 gnd
rlabel metal1 -115 -379 -115 -379 5 vdd
rlabel metal1 -148 -481 -148 -481 1 gnd
rlabel metal1 -147 -379 -147 -379 5 vdd
rlabel metal1 -374 -264 -374 -264 3 a1
rlabel metal1 -374 -476 -374 -476 3 b1
rlabel metal1 -104 -234 -104 -234 1 a1mid
rlabel metal1 -96 -445 -96 -445 1 b1mid
rlabel metal1 -353 -582 -353 -582 5 vdd
rlabel metal1 -353 -747 -353 -747 1 gnd
rlabel metal1 -301 -582 -301 -582 5 vdd
rlabel metal1 -301 -747 -301 -747 1 gnd
rlabel metal1 -249 -747 -249 -747 1 gnd
rlabel metal1 -249 -582 -249 -582 5 vdd
rlabel metal1 -197 -747 -197 -747 1 gnd
rlabel metal1 -197 -582 -197 -582 5 vdd
rlabel metal1 -121 -676 -121 -676 1 gnd
rlabel metal1 -120 -574 -120 -574 5 vdd
rlabel metal1 -153 -676 -153 -676 1 gnd
rlabel metal1 -152 -574 -152 -574 5 vdd
rlabel metal1 -354 -793 -354 -793 5 vdd
rlabel metal1 -354 -958 -354 -958 1 gnd
rlabel metal1 -302 -793 -302 -793 5 vdd
rlabel metal1 -302 -958 -302 -958 1 gnd
rlabel metal1 -250 -958 -250 -958 1 gnd
rlabel metal1 -250 -793 -250 -793 5 vdd
rlabel metal1 -198 -958 -198 -958 1 gnd
rlabel metal1 -198 -793 -198 -793 5 vdd
rlabel metal1 -122 -887 -122 -887 1 gnd
rlabel metal1 -121 -785 -121 -785 5 vdd
rlabel metal1 -154 -887 -154 -887 1 gnd
rlabel metal1 -153 -785 -153 -785 5 vdd
rlabel metal1 -380 -670 -380 -670 3 a2
rlabel metal1 -380 -882 -380 -882 3 b2
rlabel metal1 -108 -639 -108 -639 1 a2mid
rlabel metal1 -102 -851 -102 -851 1 b2mid
rlabel metal1 -140 -1487 -140 -1487 5 vdd
rlabel metal1 -141 -1589 -141 -1589 1 gnd
rlabel metal1 -108 -1487 -108 -1487 5 vdd
rlabel metal1 -109 -1589 -109 -1589 1 gnd
rlabel metal1 -185 -1495 -185 -1495 5 vdd
rlabel metal1 -185 -1660 -185 -1660 1 gnd
rlabel metal1 -237 -1495 -237 -1495 5 vdd
rlabel metal1 -237 -1660 -237 -1660 1 gnd
rlabel metal1 -289 -1660 -289 -1660 1 gnd
rlabel metal1 -289 -1495 -289 -1495 5 vdd
rlabel metal1 -341 -1660 -341 -1660 1 gnd
rlabel metal1 -341 -1495 -341 -1495 5 vdd
rlabel metal1 -139 -1276 -139 -1276 5 vdd
rlabel metal1 -140 -1378 -140 -1378 1 gnd
rlabel metal1 -107 -1276 -107 -1276 5 vdd
rlabel metal1 -108 -1378 -108 -1378 1 gnd
rlabel metal1 -184 -1284 -184 -1284 5 vdd
rlabel metal1 -184 -1449 -184 -1449 1 gnd
rlabel metal1 -236 -1284 -236 -1284 5 vdd
rlabel metal1 -236 -1449 -236 -1449 1 gnd
rlabel metal1 -288 -1449 -288 -1449 1 gnd
rlabel metal1 -288 -1284 -288 -1284 5 vdd
rlabel metal1 -340 -1449 -340 -1449 1 gnd
rlabel metal1 -340 -1284 -340 -1284 5 vdd
rlabel metal1 -98 -1342 -98 -1342 1 a3mid
rlabel metal1 -86 -1552 -86 -1552 1 b3mid
rlabel metal1 -367 -1372 -367 -1372 1 a3
rlabel metal1 -367 -1584 -367 -1584 1 b3
rlabel metal1 912 -1491 912 -1491 1 c4
rlabel metal1 1147 -1362 1147 -1362 5 vdd
rlabel metal1 1147 -1527 1147 -1527 1 gnd
rlabel metal1 1199 -1362 1199 -1362 5 vdd
rlabel metal1 1199 -1527 1199 -1527 1 gnd
rlabel metal1 1251 -1527 1251 -1527 1 gnd
rlabel metal1 1251 -1362 1251 -1362 5 vdd
rlabel metal1 1303 -1527 1303 -1527 1 gnd
rlabel metal1 1303 -1362 1303 -1362 5 vdd
rlabel metal1 1379 -1456 1379 -1456 1 gnd
rlabel metal1 1380 -1354 1380 -1354 5 vdd
rlabel metal1 1347 -1456 1347 -1456 1 gnd
rlabel metal1 1348 -1354 1348 -1354 5 vdd
rlabel metal1 1394 -1419 1394 -1419 1 cout
rlabel metal1 1393 -724 1393 -724 1 s3
rlabel metal1 1347 -658 1347 -658 5 vdd
rlabel metal1 1346 -760 1346 -760 1 gnd
rlabel metal1 1379 -658 1379 -658 5 vdd
rlabel metal1 1378 -760 1378 -760 1 gnd
rlabel metal1 1302 -666 1302 -666 5 vdd
rlabel metal1 1302 -831 1302 -831 1 gnd
rlabel metal1 1250 -666 1250 -666 5 vdd
rlabel metal1 1250 -831 1250 -831 1 gnd
rlabel metal1 1198 -831 1198 -831 1 gnd
rlabel metal1 1198 -666 1198 -666 5 vdd
rlabel metal1 1146 -831 1146 -831 1 gnd
rlabel metal1 1146 -666 1146 -666 5 vdd
rlabel metal1 1393 290 1393 290 7 s0
rlabel metal1 1349 355 1349 355 5 vdd
rlabel metal1 1348 253 1348 253 1 gnd
rlabel metal1 1381 355 1381 355 5 vdd
rlabel metal1 1380 253 1380 253 1 gnd
rlabel metal1 1304 347 1304 347 5 vdd
rlabel metal1 1304 182 1304 182 1 gnd
rlabel metal1 1252 347 1252 347 5 vdd
rlabel metal1 1252 182 1252 182 1 gnd
rlabel metal1 1200 182 1200 182 1 gnd
rlabel metal1 1200 347 1200 347 5 vdd
rlabel metal1 1148 182 1148 182 1 gnd
rlabel metal1 1148 347 1148 347 5 vdd
rlabel metal1 1392 -310 1392 -310 1 s2
rlabel metal1 1347 -244 1347 -244 5 vdd
rlabel metal1 1346 -346 1346 -346 1 gnd
rlabel metal1 1379 -244 1379 -244 5 vdd
rlabel metal1 1378 -346 1378 -346 1 gnd
rlabel metal1 1302 -252 1302 -252 5 vdd
rlabel metal1 1302 -417 1302 -417 1 gnd
rlabel metal1 1250 -252 1250 -252 5 vdd
rlabel metal1 1250 -417 1250 -417 1 gnd
rlabel metal1 1198 -417 1198 -417 1 gnd
rlabel metal1 1198 -252 1198 -252 5 vdd
rlabel metal1 1146 -417 1146 -417 1 gnd
rlabel metal1 1146 -252 1146 -252 5 vdd
rlabel metal1 893 -383 893 -383 3 vdd
rlabel metal1 995 -382 995 -382 7 gnd
rlabel metal1 995 -331 995 -331 7 gnd
rlabel metal1 893 -332 893 -332 3 vdd
rlabel metal1 1047 -309 1047 -309 5 vdd
rlabel metal1 1046 -411 1046 -411 1 gnd
rlabel metal1 1061 -375 1061 -375 1 s2mid
rlabel metal1 1060 38 1060 38 1 s1mid
rlabel metal1 1046 1 1046 1 1 gnd
rlabel metal1 1047 103 1047 103 5 vdd
rlabel metal1 893 80 893 80 3 vdd
rlabel metal1 995 81 995 81 7 gnd
rlabel metal1 995 30 995 30 7 gnd
rlabel metal1 893 29 893 29 3 vdd
rlabel metal1 893 210 893 210 3 vdd
rlabel metal1 995 211 995 211 7 gnd
rlabel metal1 995 262 995 262 7 gnd
rlabel metal1 893 261 893 261 3 vdd
rlabel metal1 1047 284 1047 284 5 vdd
rlabel metal1 1046 182 1046 182 1 gnd
rlabel metal1 1058 218 1058 218 1 s0mid
rlabel metal1 1393 89 1393 89 1 s1
rlabel metal1 1348 155 1348 155 5 vdd
rlabel metal1 1347 53 1347 53 1 gnd
rlabel metal1 1380 155 1380 155 5 vdd
rlabel metal1 1379 53 1379 53 1 gnd
rlabel metal1 1303 147 1303 147 5 vdd
rlabel metal1 1303 -18 1303 -18 1 gnd
rlabel metal1 1251 147 1251 147 5 vdd
rlabel metal1 1251 -18 1251 -18 1 gnd
rlabel metal1 1199 -18 1199 -18 1 gnd
rlabel metal1 1199 147 1199 147 5 vdd
rlabel metal1 1147 -18 1147 -18 1 gnd
rlabel metal1 1147 147 1147 147 5 vdd
rlabel metal1 1062 -807 1062 -807 1 s3mid
rlabel metal1 894 -815 894 -815 3 vdd
rlabel metal1 996 -814 996 -814 7 gnd
rlabel metal1 996 -763 996 -763 7 gnd
rlabel metal1 894 -764 894 -764 3 vdd
rlabel metal1 1048 -741 1048 -741 5 vdd
rlabel metal1 1047 -843 1047 -843 1 gnd
rlabel metal1 -95 366 -95 366 1 clk
rlabel metal1 1418 263 1418 263 1 gnd
rlabel metal1 1419 335 1419 335 5 vdd
rlabel metal1 1417 63 1417 63 1 gnd
rlabel metal1 1418 135 1418 135 5 vdd
rlabel metal1 1416 -336 1416 -336 1 gnd
rlabel metal1 1417 -264 1417 -264 5 vdd
rlabel metal1 1417 -1446 1417 -1446 1 gnd
rlabel metal1 1418 -1374 1418 -1374 5 vdd
rlabel metal1 1416 -750 1416 -750 1 gnd
rlabel metal1 1417 -678 1417 -678 5 vdd
<< end >>
